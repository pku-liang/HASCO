module MultiDimTime(
  input         clock,
  input         reset,
  input         io_in,
  output [1:0]  io_out_0,
  output [1:0]  io_out_1,
  output [17:0] io_index_0,
  output [17:0] io_index_1
);
  reg [15:0] regs_0; // @[mem.scala 68:12]
  reg [31:0] _RAND_0;
  reg [15:0] regs_1; // @[mem.scala 68:12]
  reg [31:0] _RAND_1;
  wire [15:0] _GEN_4 = {{15'd0}, io_in}; // @[mem.scala 70:42]
  wire [15:0] _T_1 = regs_0 + _GEN_4; // @[mem.scala 70:42]
  wire  back_0 = _T_1 == 16'h1; // @[mem.scala 70:48]
  wire [15:0] _T_3 = regs_1 + _GEN_4; // @[mem.scala 70:42]
  wire  back_1 = _T_3 == 16'h8; // @[mem.scala 70:48]
  wire  _T_4 = ~back_0; // @[mem.scala 77:20]
  wire [1:0] _T_5 = {_T_4, 1'h0}; // @[mem.scala 77:31]
  wire  _T_6 = ~back_1; // @[mem.scala 77:40]
  wire [1:0] _GEN_6 = {{1'd0}, _T_6}; // @[mem.scala 77:37]
  wire  _GEN_3 = back_0 ? 1'h0 : io_in; // @[mem.scala 87:16]
  assign io_out_0 = {{1'd0}, _GEN_3}; // @[mem.scala 89:15 mem.scala 92:15]
  assign io_out_1 = _T_5 | _GEN_6; // @[mem.scala 77:15]
  assign io_index_0 = {{2'd0}, regs_0}; // @[mem.scala 86:15]
  assign io_index_1 = {{2'd0}, regs_1}; // @[mem.scala 74:17]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  regs_0 = _RAND_0[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  regs_1 = _RAND_1[15:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`endif // SYNTHESIS
  always @(posedge clock) begin
    if (reset) begin
      regs_0 <= 16'h0;
    end else if (back_0) begin
      regs_0 <= 16'h0;
    end else begin
      regs_0 <= _T_1;
    end
    if (reset) begin
      regs_1 <= 16'h0;
    end else if (back_0) begin
      if (back_1) begin
        regs_1 <= 16'h0;
      end else begin
        regs_1 <= _T_3;
      end
    end
  end
endmodule
module ComputeCell_Latency(
  input        clock,
  input        reset,
  input  [7:0] io_data_2_in,
  output [7:0] io_data_2_out,
  input  [7:0] io_data_1_in,
  output [7:0] io_data_1_out,
  input  [7:0] io_data_0_in,
  output [7:0] io_data_0_out
);
  wire  _T_4 = ~reset; // @[cell.scala 111:9]
  reg [7:0] delay_a_0; // @[Reg.scala 27:20]
  reg [31:0] _RAND_0;
  reg [7:0] delay_b_0; // @[Reg.scala 27:20]
  reg [31:0] _RAND_1;
  reg [7:0] delay_c_0; // @[Reg.scala 27:20]
  reg [31:0] _RAND_2;
  wire [15:0] _T_11 = delay_a_0 * delay_b_0; // @[cell.scala 135:63]
  wire [15:0] _GEN_3 = {{8'd0}, delay_c_0}; // @[cell.scala 135:50]
  wire [15:0] _T_13 = _GEN_3 + _T_11; // @[cell.scala 135:50]
  assign io_data_2_out = io_data_2_in; // @[cell.scala 140:18]
  assign io_data_1_out = io_data_1_in; // @[cell.scala 139:18]
  assign io_data_0_out = _T_13[7:0]; // @[cell.scala 138:18]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  delay_a_0 = _RAND_0[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  delay_b_0 = _RAND_1[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  delay_c_0 = _RAND_2[7:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`endif // SYNTHESIS
  always @(posedge clock) begin
    if (reset) begin
      delay_a_0 <= 8'h0;
    end else begin
      delay_a_0 <= io_data_1_in;
    end
    if (reset) begin
      delay_b_0 <= 8'h0;
    end else begin
      delay_b_0 <= io_data_2_in;
    end
    if (reset) begin
      delay_c_0 <= 8'h0;
    end else begin
      delay_c_0 <= io_data_0_in;
    end
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_4) begin
          $fwrite(32'h80000002,"HeterogeneousBag(0 -> AnonymousBundle(in -> %d, out -> %d), 1 -> AnonymousBundle(in -> %d, out -> %d), 2 -> AnonymousBundle(in -> %d, out -> %d))\n",io_data_0_in,io_data_0_out,io_data_1_in,io_data_1_out,io_data_2_in,io_data_2_out); // @[cell.scala 111:9]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
  end
endmodule
module SystolicOutput(
  input        io_port_in_valid,
  input  [7:0] io_port_in_bits,
  output       io_port_out_valid,
  output [7:0] io_port_out_bits,
  input        io_from_cell_valid,
  input  [7:0] io_from_cell_bits,
  output       io_to_cell_valid,
  output [7:0] io_to_cell_bits
);
  assign io_port_out_valid = io_from_cell_valid; // @[pe_modules.scala 111:15]
  assign io_port_out_bits = io_from_cell_bits; // @[pe_modules.scala 111:15]
  assign io_to_cell_valid = io_port_in_valid; // @[pe_modules.scala 110:14]
  assign io_to_cell_bits = io_port_in_bits; // @[pe_modules.scala 110:14]
endmodule
module StationaryInput_Pipeline(
  input        clock,
  input        reset,
  input        io_port_in_valid,
  input  [7:0] io_port_in_bits,
  output       io_port_out_valid,
  output [7:0] io_port_out_bits,
  output [7:0] io_to_cell_bits,
  input        io_sig_stat2trans
);
  reg  trans_valid; // @[pe_modules.scala 128:22]
  reg [31:0] _RAND_0;
  reg [7:0] trans_bits; // @[pe_modules.scala 128:22]
  reg [31:0] _RAND_1;
  reg  update_valid; // @[pe_modules.scala 131:23]
  reg [31:0] _RAND_2;
  reg [7:0] update_bits_0; // @[pe_modules.scala 131:23]
  reg [31:0] _RAND_3;
  reg  stat_valid; // @[pe_modules.scala 133:21]
  reg [31:0] _RAND_4;
  reg [7:0] stat_bits_0; // @[pe_modules.scala 133:21]
  reg [31:0] _RAND_5;
  reg  reg_stat2trans_0; // @[pe_modules.scala 135:31]
  reg [31:0] _RAND_6;
  reg [3:0] write_trans_pos; // @[pe_modules.scala 137:32]
  reg [31:0] _RAND_7;
  wire  _T_4 = ~update_valid; // @[pe_modules.scala 142:26]
  wire [3:0] _GEN_5 = {{3'd0}, trans_valid}; // @[pe_modules.scala 142:60]
  wire [3:0] _T_6 = write_trans_pos + _GEN_5; // @[pe_modules.scala 142:60]
  wire  _T_7 = _T_6 == 4'h1; // @[pe_modules.scala 142:79]
  wire  _T_13 = _T_4 & trans_valid; // @[pe_modules.scala 143:24]
  wire  _T_21 = write_trans_pos == 4'h0; // @[pe_modules.scala 149:23]
  wire  _T_22 = _T_21 & trans_valid; // @[pe_modules.scala 149:45]
  wire  _GEN_1 = _T_22 | update_valid; // @[pe_modules.scala 149:60]
  reg [7:0] _T_24; // @[pe_modules.scala 163:29]
  reg [31:0] _RAND_8;
  wire  _T_26 = ~reset; // @[pe_modules.scala 165:9]
  assign io_port_out_valid = update_valid; // @[pe_modules.scala 139:21]
  assign io_port_out_bits = trans_bits; // @[pe_modules.scala 140:20]
  assign io_to_cell_bits = _T_24; // @[pe_modules.scala 163:19]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  trans_valid = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  trans_bits = _RAND_1[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  update_valid = _RAND_2[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  update_bits_0 = _RAND_3[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  stat_valid = _RAND_4[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{`RANDOM}};
  stat_bits_0 = _RAND_5[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {1{`RANDOM}};
  reg_stat2trans_0 = _RAND_6[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7 = {1{`RANDOM}};
  write_trans_pos = _RAND_7[3:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8 = {1{`RANDOM}};
  _T_24 = _RAND_8[7:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`endif // SYNTHESIS
  always @(posedge clock) begin
    if (reset) begin
      trans_valid <= 1'h0;
    end else begin
      trans_valid <= io_port_in_valid;
    end
    if (reset) begin
      trans_bits <= 8'h0;
    end else begin
      trans_bits <= io_port_in_bits;
    end
    if (reset) begin
      update_valid <= 1'h0;
    end else if (reg_stat2trans_0) begin
      update_valid <= 1'h0;
    end else begin
      update_valid <= _GEN_1;
    end
    if (reset) begin
      update_bits_0 <= 8'h0;
    end else if (_T_13) begin
      update_bits_0 <= trans_bits;
    end
    if (reset) begin
      stat_valid <= 1'h0;
    end else if (reg_stat2trans_0) begin
      stat_valid <= update_valid;
    end
    if (reset) begin
      stat_bits_0 <= 8'h0;
    end else if (reg_stat2trans_0) begin
      stat_bits_0 <= update_bits_0;
    end
    if (reset) begin
      reg_stat2trans_0 <= 1'h0;
    end else begin
      reg_stat2trans_0 <= io_sig_stat2trans;
    end
    if (reset) begin
      write_trans_pos <= 4'h0;
    end else if (_T_4) begin
      if (_T_7) begin
        write_trans_pos <= 4'h0;
      end else begin
        write_trans_pos <= _T_6;
      end
    end
    if (reset) begin
      _T_24 <= 8'h0;
    end else begin
      _T_24 <= stat_bits_0;
    end
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_26) begin
          $fwrite(32'h80000002,"sig:%d, update:Valid(valid -> %d, bits -> Vec(%d)), stat:Valid(valid -> %d, bits -> Vec(%d))\n",reg_stat2trans_0,update_valid,update_bits_0,stat_valid,stat_bits_0); // @[pe_modules.scala 165:9]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
  end
endmodule
module SystolicInput(
  input        clock,
  input        reset,
  input  [7:0] io_port_in_bits,
  output [7:0] io_port_out_bits,
  output [7:0] io_to_cell_bits
);
  reg [7:0] reg_0_bits; // @[pe_modules.scala 82:20]
  reg [31:0] _RAND_0;
  reg [7:0] to_cell_delay1_bits; // @[pe_modules.scala 83:31]
  reg [31:0] _RAND_1;
  reg [7:0] to_cell_delay2_bits; // @[pe_modules.scala 84:31]
  reg [31:0] _RAND_2;
  assign io_port_out_bits = reg_0_bits; // @[pe_modules.scala 91:15]
  assign io_to_cell_bits = to_cell_delay2_bits; // @[pe_modules.scala 92:14]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  reg_0_bits = _RAND_0[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  to_cell_delay1_bits = _RAND_1[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  to_cell_delay2_bits = _RAND_2[7:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`endif // SYNTHESIS
  always @(posedge clock) begin
    if (reset) begin
      reg_0_bits <= 8'h0;
    end else begin
      reg_0_bits <= io_port_in_bits;
    end
    if (reset) begin
      to_cell_delay1_bits <= 8'h0;
    end else begin
      to_cell_delay1_bits <= reg_0_bits;
    end
    if (reset) begin
      to_cell_delay2_bits <= 8'h0;
    end else begin
      to_cell_delay2_bits <= to_cell_delay1_bits;
    end
  end
endmodule
module PE(
  input        clock,
  input        reset,
  input  [7:0] io_data_2_in_bits,
  output [7:0] io_data_2_out_bits,
  input        io_data_1_in_valid,
  input  [7:0] io_data_1_in_bits,
  output       io_data_1_out_valid,
  output [7:0] io_data_1_out_bits,
  input        io_data_0_in_valid,
  input  [7:0] io_data_0_in_bits,
  output       io_data_0_out_valid,
  output [7:0] io_data_0_out_bits,
  input        io_sig_stat2trans
);
  wire  ComputeCell_Latency_clock; // @[pe.scala 37:18]
  wire  ComputeCell_Latency_reset; // @[pe.scala 37:18]
  wire [7:0] ComputeCell_Latency_io_data_2_in; // @[pe.scala 37:18]
  wire [7:0] ComputeCell_Latency_io_data_2_out; // @[pe.scala 37:18]
  wire [7:0] ComputeCell_Latency_io_data_1_in; // @[pe.scala 37:18]
  wire [7:0] ComputeCell_Latency_io_data_1_out; // @[pe.scala 37:18]
  wire [7:0] ComputeCell_Latency_io_data_0_in; // @[pe.scala 37:18]
  wire [7:0] ComputeCell_Latency_io_data_0_out; // @[pe.scala 37:18]
  wire  SystolicOutput_io_port_in_valid; // @[pe.scala 39:11]
  wire [7:0] SystolicOutput_io_port_in_bits; // @[pe.scala 39:11]
  wire  SystolicOutput_io_port_out_valid; // @[pe.scala 39:11]
  wire [7:0] SystolicOutput_io_port_out_bits; // @[pe.scala 39:11]
  wire  SystolicOutput_io_from_cell_valid; // @[pe.scala 39:11]
  wire [7:0] SystolicOutput_io_from_cell_bits; // @[pe.scala 39:11]
  wire  SystolicOutput_io_to_cell_valid; // @[pe.scala 39:11]
  wire [7:0] SystolicOutput_io_to_cell_bits; // @[pe.scala 39:11]
  wire  StationaryInput_Pipeline_clock; // @[pe.scala 39:11]
  wire  StationaryInput_Pipeline_reset; // @[pe.scala 39:11]
  wire  StationaryInput_Pipeline_io_port_in_valid; // @[pe.scala 39:11]
  wire [7:0] StationaryInput_Pipeline_io_port_in_bits; // @[pe.scala 39:11]
  wire  StationaryInput_Pipeline_io_port_out_valid; // @[pe.scala 39:11]
  wire [7:0] StationaryInput_Pipeline_io_port_out_bits; // @[pe.scala 39:11]
  wire [7:0] StationaryInput_Pipeline_io_to_cell_bits; // @[pe.scala 39:11]
  wire  StationaryInput_Pipeline_io_sig_stat2trans; // @[pe.scala 39:11]
  wire  SystolicInput_clock; // @[pe.scala 39:11]
  wire  SystolicInput_reset; // @[pe.scala 39:11]
  wire [7:0] SystolicInput_io_port_in_bits; // @[pe.scala 39:11]
  wire [7:0] SystolicInput_io_port_out_bits; // @[pe.scala 39:11]
  wire [7:0] SystolicInput_io_to_cell_bits; // @[pe.scala 39:11]
  wire  _T_4 = ~reset; // @[pe.scala 28:9]
  reg  _T_5; // @[Reg.scala 15:16]
  reg [31:0] _RAND_0;
  ComputeCell_Latency ComputeCell_Latency ( // @[pe.scala 37:18]
    .clock(ComputeCell_Latency_clock),
    .reset(ComputeCell_Latency_reset),
    .io_data_2_in(ComputeCell_Latency_io_data_2_in),
    .io_data_2_out(ComputeCell_Latency_io_data_2_out),
    .io_data_1_in(ComputeCell_Latency_io_data_1_in),
    .io_data_1_out(ComputeCell_Latency_io_data_1_out),
    .io_data_0_in(ComputeCell_Latency_io_data_0_in),
    .io_data_0_out(ComputeCell_Latency_io_data_0_out)
  );
  SystolicOutput SystolicOutput ( // @[pe.scala 39:11]
    .io_port_in_valid(SystolicOutput_io_port_in_valid),
    .io_port_in_bits(SystolicOutput_io_port_in_bits),
    .io_port_out_valid(SystolicOutput_io_port_out_valid),
    .io_port_out_bits(SystolicOutput_io_port_out_bits),
    .io_from_cell_valid(SystolicOutput_io_from_cell_valid),
    .io_from_cell_bits(SystolicOutput_io_from_cell_bits),
    .io_to_cell_valid(SystolicOutput_io_to_cell_valid),
    .io_to_cell_bits(SystolicOutput_io_to_cell_bits)
  );
  StationaryInput_Pipeline StationaryInput_Pipeline ( // @[pe.scala 39:11]
    .clock(StationaryInput_Pipeline_clock),
    .reset(StationaryInput_Pipeline_reset),
    .io_port_in_valid(StationaryInput_Pipeline_io_port_in_valid),
    .io_port_in_bits(StationaryInput_Pipeline_io_port_in_bits),
    .io_port_out_valid(StationaryInput_Pipeline_io_port_out_valid),
    .io_port_out_bits(StationaryInput_Pipeline_io_port_out_bits),
    .io_to_cell_bits(StationaryInput_Pipeline_io_to_cell_bits),
    .io_sig_stat2trans(StationaryInput_Pipeline_io_sig_stat2trans)
  );
  SystolicInput SystolicInput ( // @[pe.scala 39:11]
    .clock(SystolicInput_clock),
    .reset(SystolicInput_reset),
    .io_port_in_bits(SystolicInput_io_port_in_bits),
    .io_port_out_bits(SystolicInput_io_port_out_bits),
    .io_to_cell_bits(SystolicInput_io_to_cell_bits)
  );
  assign io_data_2_out_bits = SystolicInput_io_port_out_bits; // @[pe.scala 42:17]
  assign io_data_1_out_valid = StationaryInput_Pipeline_io_port_out_valid; // @[pe.scala 42:17]
  assign io_data_1_out_bits = StationaryInput_Pipeline_io_port_out_bits; // @[pe.scala 42:17]
  assign io_data_0_out_valid = SystolicOutput_io_port_out_valid; // @[pe.scala 42:17]
  assign io_data_0_out_bits = SystolicOutput_io_port_out_bits; // @[pe.scala 42:17]
  assign ComputeCell_Latency_clock = clock;
  assign ComputeCell_Latency_reset = reset;
  assign ComputeCell_Latency_io_data_2_in = SystolicInput_io_to_cell_bits; // @[pe.scala 43:19]
  assign ComputeCell_Latency_io_data_1_in = StationaryInput_Pipeline_io_to_cell_bits; // @[pe.scala 43:19]
  assign ComputeCell_Latency_io_data_0_in = SystolicOutput_io_to_cell_bits; // @[pe.scala 43:19]
  assign SystolicOutput_io_port_in_valid = io_data_0_in_valid; // @[pe.scala 42:17]
  assign SystolicOutput_io_port_in_bits = io_data_0_in_bits; // @[pe.scala 42:17]
  assign SystolicOutput_io_from_cell_valid = _T_5; // @[pe.scala 46:34]
  assign SystolicOutput_io_from_cell_bits = ComputeCell_Latency_io_data_0_out; // @[pe.scala 45:33]
  assign StationaryInput_Pipeline_clock = clock;
  assign StationaryInput_Pipeline_reset = reset;
  assign StationaryInput_Pipeline_io_port_in_valid = io_data_1_in_valid; // @[pe.scala 42:17]
  assign StationaryInput_Pipeline_io_port_in_bits = io_data_1_in_bits; // @[pe.scala 42:17]
  assign StationaryInput_Pipeline_io_sig_stat2trans = io_sig_stat2trans; // @[pe.scala 50:33]
  assign SystolicInput_clock = clock;
  assign SystolicInput_reset = reset;
  assign SystolicInput_io_port_in_bits = io_data_2_in_bits; // @[pe.scala 42:17]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _T_5 = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`endif // SYNTHESIS
  always @(posedge clock) begin
    _T_5 <= SystolicOutput_io_to_cell_valid;
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_4) begin
          $fwrite(32'h80000002,"data0=%d,data1=%d,data2=%d,sig=%d\n",io_data_0_in_bits,io_data_1_in_bits,io_data_2_in_bits,io_sig_stat2trans); // @[pe.scala 28:9]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
  end
endmodule
module PENetwork(
  input        io_to_pes_0_out_valid,
  input  [7:0] io_to_pes_0_out_bits,
  output       io_to_pes_1_in_valid,
  output [7:0] io_to_pes_1_in_bits,
  input        io_to_pes_1_out_valid,
  input  [7:0] io_to_pes_1_out_bits,
  output       io_to_pes_2_in_valid,
  output [7:0] io_to_pes_2_in_bits,
  input        io_to_pes_2_out_valid,
  input  [7:0] io_to_pes_2_out_bits,
  output       io_to_pes_3_in_valid,
  output [7:0] io_to_pes_3_in_bits,
  input        io_to_pes_3_out_valid,
  input  [7:0] io_to_pes_3_out_bits,
  output       io_to_pes_4_in_valid,
  output [7:0] io_to_pes_4_in_bits,
  input        io_to_pes_4_out_valid,
  input  [7:0] io_to_pes_4_out_bits,
  output       io_to_pes_5_in_valid,
  output [7:0] io_to_pes_5_in_bits,
  input        io_to_pes_5_out_valid,
  input  [7:0] io_to_pes_5_out_bits,
  output       io_to_pes_6_in_valid,
  output [7:0] io_to_pes_6_in_bits,
  input        io_to_pes_6_out_valid,
  input  [7:0] io_to_pes_6_out_bits,
  output       io_to_pes_7_in_valid,
  output [7:0] io_to_pes_7_in_bits,
  input        io_to_pes_7_out_valid,
  input  [7:0] io_to_pes_7_out_bits,
  output       io_to_mem_valid,
  output [7:0] io_to_mem_bits
);
  assign io_to_pes_1_in_valid = io_to_pes_0_out_valid; // @[pearray.scala 38:23]
  assign io_to_pes_1_in_bits = io_to_pes_0_out_bits; // @[pearray.scala 38:23]
  assign io_to_pes_2_in_valid = io_to_pes_1_out_valid; // @[pearray.scala 38:23]
  assign io_to_pes_2_in_bits = io_to_pes_1_out_bits; // @[pearray.scala 38:23]
  assign io_to_pes_3_in_valid = io_to_pes_2_out_valid; // @[pearray.scala 38:23]
  assign io_to_pes_3_in_bits = io_to_pes_2_out_bits; // @[pearray.scala 38:23]
  assign io_to_pes_4_in_valid = io_to_pes_3_out_valid; // @[pearray.scala 38:23]
  assign io_to_pes_4_in_bits = io_to_pes_3_out_bits; // @[pearray.scala 38:23]
  assign io_to_pes_5_in_valid = io_to_pes_4_out_valid; // @[pearray.scala 38:23]
  assign io_to_pes_5_in_bits = io_to_pes_4_out_bits; // @[pearray.scala 38:23]
  assign io_to_pes_6_in_valid = io_to_pes_5_out_valid; // @[pearray.scala 38:23]
  assign io_to_pes_6_in_bits = io_to_pes_5_out_bits; // @[pearray.scala 38:23]
  assign io_to_pes_7_in_valid = io_to_pes_6_out_valid; // @[pearray.scala 38:23]
  assign io_to_pes_7_in_bits = io_to_pes_6_out_bits; // @[pearray.scala 38:23]
  assign io_to_mem_valid = io_to_pes_7_out_valid; // @[pearray.scala 45:17]
  assign io_to_mem_bits = io_to_pes_7_out_bits; // @[pearray.scala 45:17]
endmodule
module PENetwork_16(
  output       io_to_pes_0_in_valid,
  output [7:0] io_to_pes_0_in_bits,
  input        io_to_pes_0_out_valid,
  input  [7:0] io_to_pes_0_out_bits,
  output       io_to_pes_1_in_valid,
  output [7:0] io_to_pes_1_in_bits,
  input        io_to_pes_1_out_valid,
  input  [7:0] io_to_pes_1_out_bits,
  output       io_to_pes_2_in_valid,
  output [7:0] io_to_pes_2_in_bits,
  input        io_to_pes_2_out_valid,
  input  [7:0] io_to_pes_2_out_bits,
  output       io_to_pes_3_in_valid,
  output [7:0] io_to_pes_3_in_bits,
  input        io_to_pes_3_out_valid,
  input  [7:0] io_to_pes_3_out_bits,
  output       io_to_pes_4_in_valid,
  output [7:0] io_to_pes_4_in_bits,
  input        io_to_pes_4_out_valid,
  input  [7:0] io_to_pes_4_out_bits,
  output       io_to_pes_5_in_valid,
  output [7:0] io_to_pes_5_in_bits,
  input        io_to_pes_5_out_valid,
  input  [7:0] io_to_pes_5_out_bits,
  output       io_to_pes_6_in_valid,
  output [7:0] io_to_pes_6_in_bits,
  input        io_to_pes_6_out_valid,
  input  [7:0] io_to_pes_6_out_bits,
  output       io_to_pes_7_in_valid,
  output [7:0] io_to_pes_7_in_bits,
  input        io_to_mem_valid,
  input  [7:0] io_to_mem_bits
);
  assign io_to_pes_0_in_valid = io_to_mem_valid; // @[pearray.scala 41:23]
  assign io_to_pes_0_in_bits = io_to_mem_bits; // @[pearray.scala 41:23]
  assign io_to_pes_1_in_valid = io_to_pes_0_out_valid; // @[pearray.scala 38:23]
  assign io_to_pes_1_in_bits = io_to_pes_0_out_bits; // @[pearray.scala 38:23]
  assign io_to_pes_2_in_valid = io_to_pes_1_out_valid; // @[pearray.scala 38:23]
  assign io_to_pes_2_in_bits = io_to_pes_1_out_bits; // @[pearray.scala 38:23]
  assign io_to_pes_3_in_valid = io_to_pes_2_out_valid; // @[pearray.scala 38:23]
  assign io_to_pes_3_in_bits = io_to_pes_2_out_bits; // @[pearray.scala 38:23]
  assign io_to_pes_4_in_valid = io_to_pes_3_out_valid; // @[pearray.scala 38:23]
  assign io_to_pes_4_in_bits = io_to_pes_3_out_bits; // @[pearray.scala 38:23]
  assign io_to_pes_5_in_valid = io_to_pes_4_out_valid; // @[pearray.scala 38:23]
  assign io_to_pes_5_in_bits = io_to_pes_4_out_bits; // @[pearray.scala 38:23]
  assign io_to_pes_6_in_valid = io_to_pes_5_out_valid; // @[pearray.scala 38:23]
  assign io_to_pes_6_in_bits = io_to_pes_5_out_bits; // @[pearray.scala 38:23]
  assign io_to_pes_7_in_valid = io_to_pes_6_out_valid; // @[pearray.scala 38:23]
  assign io_to_pes_7_in_bits = io_to_pes_6_out_bits; // @[pearray.scala 38:23]
endmodule
module PENetwork_32(
  output [7:0] io_to_pes_0_in_bits,
  input  [7:0] io_to_pes_0_out_bits,
  output [7:0] io_to_pes_1_in_bits,
  input  [7:0] io_to_pes_1_out_bits,
  output [7:0] io_to_pes_2_in_bits,
  input  [7:0] io_to_pes_2_out_bits,
  output [7:0] io_to_pes_3_in_bits,
  input  [7:0] io_to_pes_3_out_bits,
  output [7:0] io_to_pes_4_in_bits,
  input  [7:0] io_to_pes_4_out_bits,
  output [7:0] io_to_pes_5_in_bits,
  input  [7:0] io_to_pes_5_out_bits,
  output [7:0] io_to_pes_6_in_bits,
  input  [7:0] io_to_pes_6_out_bits,
  output [7:0] io_to_pes_7_in_bits,
  input  [7:0] io_to_pes_7_out_bits,
  output [7:0] io_to_pes_8_in_bits,
  input  [7:0] io_to_pes_8_out_bits,
  output [7:0] io_to_pes_9_in_bits,
  input  [7:0] io_to_pes_9_out_bits,
  output [7:0] io_to_pes_10_in_bits,
  input  [7:0] io_to_pes_10_out_bits,
  output [7:0] io_to_pes_11_in_bits,
  input  [7:0] io_to_pes_11_out_bits,
  output [7:0] io_to_pes_12_in_bits,
  input  [7:0] io_to_pes_12_out_bits,
  output [7:0] io_to_pes_13_in_bits,
  input  [7:0] io_to_pes_13_out_bits,
  output [7:0] io_to_pes_14_in_bits,
  input  [7:0] io_to_pes_14_out_bits,
  output [7:0] io_to_pes_15_in_bits,
  input  [7:0] io_to_mem_bits
);
  assign io_to_pes_0_in_bits = io_to_mem_bits; // @[pearray.scala 41:23]
  assign io_to_pes_1_in_bits = io_to_pes_0_out_bits; // @[pearray.scala 38:23]
  assign io_to_pes_2_in_bits = io_to_pes_1_out_bits; // @[pearray.scala 38:23]
  assign io_to_pes_3_in_bits = io_to_pes_2_out_bits; // @[pearray.scala 38:23]
  assign io_to_pes_4_in_bits = io_to_pes_3_out_bits; // @[pearray.scala 38:23]
  assign io_to_pes_5_in_bits = io_to_pes_4_out_bits; // @[pearray.scala 38:23]
  assign io_to_pes_6_in_bits = io_to_pes_5_out_bits; // @[pearray.scala 38:23]
  assign io_to_pes_7_in_bits = io_to_pes_6_out_bits; // @[pearray.scala 38:23]
  assign io_to_pes_8_in_bits = io_to_pes_7_out_bits; // @[pearray.scala 38:23]
  assign io_to_pes_9_in_bits = io_to_pes_8_out_bits; // @[pearray.scala 38:23]
  assign io_to_pes_10_in_bits = io_to_pes_9_out_bits; // @[pearray.scala 38:23]
  assign io_to_pes_11_in_bits = io_to_pes_10_out_bits; // @[pearray.scala 38:23]
  assign io_to_pes_12_in_bits = io_to_pes_11_out_bits; // @[pearray.scala 38:23]
  assign io_to_pes_13_in_bits = io_to_pes_12_out_bits; // @[pearray.scala 38:23]
  assign io_to_pes_14_in_bits = io_to_pes_13_out_bits; // @[pearray.scala 38:23]
  assign io_to_pes_15_in_bits = io_to_pes_14_out_bits; // @[pearray.scala 38:23]
endmodule
module MultiDimMem(
  input        clock,
  input        reset,
  input        io_rd_addr_valid,
  input  [1:0] io_rd_addr_bits_0,
  input  [1:0] io_rd_addr_bits_1,
  output       io_rd_data_valid,
  output [7:0] io_rd_data_bits,
  input  [1:0] io_wr_addr_bits_0,
  input  [1:0] io_wr_addr_bits_1,
  input        io_wr_data_valid,
  input  [7:0] io_wr_data_bits
);
  reg [8:0] mem [0:7]; // @[mem.scala 106:24]
  reg [31:0] _RAND_0;
  wire [8:0] mem_mem_output_data; // @[mem.scala 106:24]
  wire [2:0] mem_mem_output_addr; // @[mem.scala 106:24]
  wire [8:0] mem__T_43_data; // @[mem.scala 106:24]
  wire [2:0] mem__T_43_addr; // @[mem.scala 106:24]
  wire  mem__T_43_mask; // @[mem.scala 106:24]
  wire  mem__T_43_en; // @[mem.scala 106:24]
  reg  mem_mem_output_en_pipe_0;
  reg [31:0] _RAND_1;
  reg [2:0] mem_mem_output_addr_pipe_0;
  reg [31:0] _RAND_2;
  reg  rd_addr_reg_valid; // @[mem.scala 107:28]
  reg [31:0] _RAND_3;
  reg [15:0] rd_addr_reg_bits_1; // @[mem.scala 107:28]
  reg [31:0] _RAND_4;
  reg [15:0] rd_addr_reg_bits_0; // @[mem.scala 107:28]
  reg [31:0] _RAND_5;
  wire [15:0] _T_6 = rd_addr_reg_bits_0 + 16'h1; // @[mem.scala 118:102]
  wire  _T_7 = 2'h1 == io_rd_addr_bits_0; // @[Mux.scala 68:19]
  wire  _T_9 = 2'h0 == io_rd_addr_bits_0; // @[Mux.scala 68:19]
  wire [15:0] _T_11 = rd_addr_reg_bits_1 + 16'h1; // @[mem.scala 118:102]
  wire  _T_12 = 2'h1 == io_rd_addr_bits_1; // @[Mux.scala 68:19]
  wire  _T_14 = 2'h0 == io_rd_addr_bits_1; // @[Mux.scala 68:19]
  wire [15:0] mem_rd_addr = rd_addr_reg_bits_0 + rd_addr_reg_bits_1; // @[mem.scala 122:46]
  reg  mem_req_valid; // @[mem.scala 129:30]
  reg [31:0] _RAND_6;
  reg [15:0] wr_addr_reg_bits_1; // @[mem.scala 131:28]
  reg [31:0] _RAND_7;
  reg [15:0] wr_addr_reg_bits_0; // @[mem.scala 131:28]
  reg [31:0] _RAND_8;
  wire [15:0] _T_22 = wr_addr_reg_bits_0 + 16'h1; // @[mem.scala 143:102]
  wire  _T_23 = 2'h1 == io_wr_addr_bits_0; // @[Mux.scala 68:19]
  wire  _T_25 = 2'h0 == io_wr_addr_bits_0; // @[Mux.scala 68:19]
  wire [15:0] _T_27 = wr_addr_reg_bits_1 + 16'h1; // @[mem.scala 143:102]
  wire  _T_28 = 2'h1 == io_wr_addr_bits_1; // @[Mux.scala 68:19]
  wire  _T_30 = 2'h0 == io_wr_addr_bits_1; // @[Mux.scala 68:19]
  wire [15:0] mem_wr_addr = wr_addr_reg_bits_0 + wr_addr_reg_bits_1; // @[mem.scala 147:46]
  reg  wr_data_1_valid; // @[mem.scala 156:26]
  reg [31:0] _RAND_9;
  reg [7:0] wr_data_1_bits; // @[mem.scala 156:26]
  reg [31:0] _RAND_10;
  reg  wr_data_2_valid; // @[mem.scala 163:26]
  reg [31:0] _RAND_11;
  reg [7:0] wr_data_2_bits; // @[mem.scala 163:26]
  reg [31:0] _RAND_12;
  reg [15:0] wr_addr_2; // @[mem.scala 165:26]
  reg [31:0] _RAND_13;
  reg [7:0] wr_data_final; // @[mem.scala 174:30]
  reg [31:0] _RAND_14;
  reg [15:0] wr_addr_3; // @[mem.scala 175:26]
  reg [31:0] _RAND_15;
  reg  wr_valid_3; // @[mem.scala 176:27]
  reg [31:0] _RAND_16;
  wire [8:0] _GEN_9 = {wr_valid_3, 8'h0}; // @[mem.scala 181:38]
  wire [15:0] _T_39 = {{7'd0}, _GEN_9}; // @[mem.scala 181:38]
  wire [15:0] _GEN_10 = {{8'd0}, wr_data_final}; // @[mem.scala 181:52]
  wire [15:0] _T_40 = _T_39 | _GEN_10; // @[mem.scala 181:52]
  reg  _T_46; // @[mem.scala 186:30]
  reg [31:0] _RAND_17;
  reg [7:0] _T_49; // @[mem.scala 187:29]
  reg [31:0] _RAND_18;
  wire  _T_51 = ~reset; // @[mem.scala 191:9]
  assign mem_mem_output_addr = mem_mem_output_addr_pipe_0;
  assign mem_mem_output_data = mem[mem_mem_output_addr]; // @[mem.scala 106:24]
  assign mem__T_43_data = _T_40[8:0];
  assign mem__T_43_addr = wr_addr_3[2:0];
  assign mem__T_43_mask = 1'h1;
  assign mem__T_43_en = wr_valid_3;
  assign io_rd_data_valid = _T_46; // @[mem.scala 186:20]
  assign io_rd_data_bits = _T_49; // @[mem.scala 187:19]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  _RAND_0 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 8; initvar = initvar+1)
    mem[initvar] = _RAND_0[8:0];
  `endif // RANDOMIZE_MEM_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  mem_mem_output_en_pipe_0 = _RAND_1[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  mem_mem_output_addr_pipe_0 = _RAND_2[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  rd_addr_reg_valid = _RAND_3[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  rd_addr_reg_bits_1 = _RAND_4[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{`RANDOM}};
  rd_addr_reg_bits_0 = _RAND_5[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {1{`RANDOM}};
  mem_req_valid = _RAND_6[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7 = {1{`RANDOM}};
  wr_addr_reg_bits_1 = _RAND_7[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8 = {1{`RANDOM}};
  wr_addr_reg_bits_0 = _RAND_8[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9 = {1{`RANDOM}};
  wr_data_1_valid = _RAND_9[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10 = {1{`RANDOM}};
  wr_data_1_bits = _RAND_10[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11 = {1{`RANDOM}};
  wr_data_2_valid = _RAND_11[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_12 = {1{`RANDOM}};
  wr_data_2_bits = _RAND_12[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_13 = {1{`RANDOM}};
  wr_addr_2 = _RAND_13[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_14 = {1{`RANDOM}};
  wr_data_final = _RAND_14[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_15 = {1{`RANDOM}};
  wr_addr_3 = _RAND_15[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_16 = {1{`RANDOM}};
  wr_valid_3 = _RAND_16[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_17 = {1{`RANDOM}};
  _T_46 = _RAND_17[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_18 = {1{`RANDOM}};
  _T_49 = _RAND_18[7:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`endif // SYNTHESIS
  always @(posedge clock) begin
    if(mem__T_43_en & mem__T_43_mask) begin
      mem[mem__T_43_addr] <= mem__T_43_data; // @[mem.scala 106:24]
    end
    mem_mem_output_en_pipe_0 <= rd_addr_reg_valid;
    if (rd_addr_reg_valid) begin
      mem_mem_output_addr_pipe_0 <= mem_rd_addr[2:0];
    end
    if (reset) begin
      rd_addr_reg_valid <= 1'h0;
    end else begin
      rd_addr_reg_valid <= io_rd_addr_valid;
    end
    if (reset) begin
      rd_addr_reg_bits_1 <= 16'h0;
    end else if (_T_14) begin
      rd_addr_reg_bits_1 <= 16'h0;
    end else if (_T_12) begin
      rd_addr_reg_bits_1 <= _T_11;
    end
    if (reset) begin
      rd_addr_reg_bits_0 <= 16'h0;
    end else if (_T_9) begin
      rd_addr_reg_bits_0 <= 16'h0;
    end else if (_T_7) begin
      rd_addr_reg_bits_0 <= _T_6;
    end
    if (reset) begin
      mem_req_valid <= 1'h0;
    end else begin
      mem_req_valid <= rd_addr_reg_valid;
    end
    if (reset) begin
      wr_addr_reg_bits_1 <= 16'h0;
    end else if (_T_30) begin
      wr_addr_reg_bits_1 <= 16'h0;
    end else if (_T_28) begin
      wr_addr_reg_bits_1 <= _T_27;
    end
    if (reset) begin
      wr_addr_reg_bits_0 <= 16'h0;
    end else if (_T_25) begin
      wr_addr_reg_bits_0 <= 16'h0;
    end else if (_T_23) begin
      wr_addr_reg_bits_0 <= _T_22;
    end
    if (reset) begin
      wr_data_1_valid <= 1'h0;
    end else begin
      wr_data_1_valid <= io_wr_data_valid;
    end
    if (reset) begin
      wr_data_1_bits <= 8'h0;
    end else begin
      wr_data_1_bits <= io_wr_data_bits;
    end
    if (reset) begin
      wr_data_2_valid <= 1'h0;
    end else begin
      wr_data_2_valid <= wr_data_1_valid;
    end
    if (reset) begin
      wr_data_2_bits <= 8'h0;
    end else begin
      wr_data_2_bits <= wr_data_1_bits;
    end
    if (reset) begin
      wr_addr_2 <= 16'h0;
    end else begin
      wr_addr_2 <= mem_wr_addr;
    end
    wr_data_final <= wr_data_2_bits;
    if (reset) begin
      wr_addr_3 <= 16'h0;
    end else begin
      wr_addr_3 <= wr_addr_2;
    end
    wr_valid_3 <= wr_data_2_valid;
    _T_46 <= mem_req_valid & mem_mem_output_data[8];
    if (mem_req_valid) begin
      _T_49 <= mem_mem_output_data[7:0];
    end else begin
      _T_49 <= 8'h0;
    end
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_51) begin
          $fwrite(32'h80000002,"io.rd_addr: %d %d, rd_addr: %d, rd_data: %d %d\n",io_rd_addr_bits_0,io_rd_addr_bits_1,mem_rd_addr,io_rd_data_valid,io_rd_data_bits); // @[mem.scala 191:9]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_51) begin
          $fwrite(32'h80000002,"wr_addr: %d, wr_addr: %d %d\n",wr_addr_3,wr_data_final,wr_valid_3); // @[mem.scala 192:9]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
  end
endmodule
module MemController(
  input        clock,
  input        reset,
  input        io_rd_valid,
  input        io_wr_valid,
  output       io_rd_data_valid,
  output [7:0] io_rd_data_bits,
  input        io_wr_data_valid,
  input  [7:0] io_wr_data_bits
);
  wire  MultiDimMem_clock; // @[mem.scala 33:19]
  wire  MultiDimMem_reset; // @[mem.scala 33:19]
  wire  MultiDimMem_io_rd_addr_valid; // @[mem.scala 33:19]
  wire [1:0] MultiDimMem_io_rd_addr_bits_0; // @[mem.scala 33:19]
  wire [1:0] MultiDimMem_io_rd_addr_bits_1; // @[mem.scala 33:19]
  wire  MultiDimMem_io_rd_data_valid; // @[mem.scala 33:19]
  wire [7:0] MultiDimMem_io_rd_data_bits; // @[mem.scala 33:19]
  wire [1:0] MultiDimMem_io_wr_addr_bits_0; // @[mem.scala 33:19]
  wire [1:0] MultiDimMem_io_wr_addr_bits_1; // @[mem.scala 33:19]
  wire  MultiDimMem_io_wr_data_valid; // @[mem.scala 33:19]
  wire [7:0] MultiDimMem_io_wr_data_bits; // @[mem.scala 33:19]
  wire  MultiDimTime_clock; // @[mem.scala 34:23]
  wire  MultiDimTime_reset; // @[mem.scala 34:23]
  wire  MultiDimTime_io_in; // @[mem.scala 34:23]
  wire [1:0] MultiDimTime_io_out_0; // @[mem.scala 34:23]
  wire [1:0] MultiDimTime_io_out_1; // @[mem.scala 34:23]
  wire [17:0] MultiDimTime_io_index_0; // @[mem.scala 34:23]
  wire [17:0] MultiDimTime_io_index_1; // @[mem.scala 34:23]
  wire  MultiDimTime_1_clock; // @[mem.scala 35:23]
  wire  MultiDimTime_1_reset; // @[mem.scala 35:23]
  wire  MultiDimTime_1_io_in; // @[mem.scala 35:23]
  wire [1:0] MultiDimTime_1_io_out_0; // @[mem.scala 35:23]
  wire [1:0] MultiDimTime_1_io_out_1; // @[mem.scala 35:23]
  wire [17:0] MultiDimTime_1_io_index_0; // @[mem.scala 35:23]
  wire [17:0] MultiDimTime_1_io_index_1; // @[mem.scala 35:23]
  MultiDimMem MultiDimMem ( // @[mem.scala 33:19]
    .clock(MultiDimMem_clock),
    .reset(MultiDimMem_reset),
    .io_rd_addr_valid(MultiDimMem_io_rd_addr_valid),
    .io_rd_addr_bits_0(MultiDimMem_io_rd_addr_bits_0),
    .io_rd_addr_bits_1(MultiDimMem_io_rd_addr_bits_1),
    .io_rd_data_valid(MultiDimMem_io_rd_data_valid),
    .io_rd_data_bits(MultiDimMem_io_rd_data_bits),
    .io_wr_addr_bits_0(MultiDimMem_io_wr_addr_bits_0),
    .io_wr_addr_bits_1(MultiDimMem_io_wr_addr_bits_1),
    .io_wr_data_valid(MultiDimMem_io_wr_data_valid),
    .io_wr_data_bits(MultiDimMem_io_wr_data_bits)
  );
  MultiDimTime MultiDimTime ( // @[mem.scala 34:23]
    .clock(MultiDimTime_clock),
    .reset(MultiDimTime_reset),
    .io_in(MultiDimTime_io_in),
    .io_out_0(MultiDimTime_io_out_0),
    .io_out_1(MultiDimTime_io_out_1),
    .io_index_0(MultiDimTime_io_index_0),
    .io_index_1(MultiDimTime_io_index_1)
  );
  MultiDimTime MultiDimTime_1 ( // @[mem.scala 35:23]
    .clock(MultiDimTime_1_clock),
    .reset(MultiDimTime_1_reset),
    .io_in(MultiDimTime_1_io_in),
    .io_out_0(MultiDimTime_1_io_out_0),
    .io_out_1(MultiDimTime_1_io_out_1),
    .io_index_0(MultiDimTime_1_io_index_0),
    .io_index_1(MultiDimTime_1_io_index_1)
  );
  assign io_rd_data_valid = MultiDimMem_io_rd_data_valid; // @[mem.scala 53:14]
  assign io_rd_data_bits = MultiDimMem_io_rd_data_bits; // @[mem.scala 53:14]
  assign MultiDimMem_clock = clock;
  assign MultiDimMem_reset = reset;
  assign MultiDimMem_io_rd_addr_valid = io_rd_valid; // @[mem.scala 50:21]
  assign MultiDimMem_io_rd_addr_bits_0 = MultiDimTime_1_io_out_0; // @[mem.scala 49:20]
  assign MultiDimMem_io_rd_addr_bits_1 = MultiDimTime_1_io_out_1; // @[mem.scala 49:20]
  assign MultiDimMem_io_wr_addr_bits_0 = MultiDimTime_io_out_0; // @[mem.scala 45:20]
  assign MultiDimMem_io_wr_addr_bits_1 = MultiDimTime_io_out_1; // @[mem.scala 45:20]
  assign MultiDimMem_io_wr_data_valid = io_wr_data_valid; // @[mem.scala 54:15]
  assign MultiDimMem_io_wr_data_bits = io_wr_data_bits; // @[mem.scala 54:15]
  assign MultiDimTime_clock = clock;
  assign MultiDimTime_reset = reset;
  assign MultiDimTime_io_in = io_wr_valid; // @[mem.scala 44:14]
  assign MultiDimTime_1_clock = clock;
  assign MultiDimTime_1_reset = reset;
  assign MultiDimTime_1_io_in = io_rd_valid; // @[mem.scala 48:14]
endmodule
module PEArray(
  input        clock,
  input        reset,
  input        io_data_2_in_0_valid,
  input        io_data_2_in_0_bits_valid,
  input  [7:0] io_data_2_in_0_bits_bits,
  input        io_data_2_in_1_valid,
  input        io_data_2_in_1_bits_valid,
  input  [7:0] io_data_2_in_1_bits_bits,
  input        io_data_2_in_2_valid,
  input        io_data_2_in_2_bits_valid,
  input  [7:0] io_data_2_in_2_bits_bits,
  input        io_data_2_in_3_valid,
  input        io_data_2_in_3_bits_valid,
  input  [7:0] io_data_2_in_3_bits_bits,
  input        io_data_2_in_4_valid,
  input        io_data_2_in_4_bits_valid,
  input  [7:0] io_data_2_in_4_bits_bits,
  input        io_data_2_in_5_valid,
  input        io_data_2_in_5_bits_valid,
  input  [7:0] io_data_2_in_5_bits_bits,
  input        io_data_2_in_6_valid,
  input        io_data_2_in_6_bits_valid,
  input  [7:0] io_data_2_in_6_bits_bits,
  input        io_data_2_in_7_valid,
  input        io_data_2_in_7_bits_valid,
  input  [7:0] io_data_2_in_7_bits_bits,
  input        io_data_1_in_0_valid,
  input        io_data_1_in_0_bits_valid,
  input  [7:0] io_data_1_in_0_bits_bits,
  input        io_data_1_in_1_valid,
  input        io_data_1_in_1_bits_valid,
  input  [7:0] io_data_1_in_1_bits_bits,
  input        io_data_1_in_2_valid,
  input        io_data_1_in_2_bits_valid,
  input  [7:0] io_data_1_in_2_bits_bits,
  input        io_data_1_in_3_valid,
  input        io_data_1_in_3_bits_valid,
  input  [7:0] io_data_1_in_3_bits_bits,
  input        io_data_1_in_4_valid,
  input        io_data_1_in_4_bits_valid,
  input  [7:0] io_data_1_in_4_bits_bits,
  input        io_data_1_in_5_valid,
  input        io_data_1_in_5_bits_valid,
  input  [7:0] io_data_1_in_5_bits_bits,
  input        io_data_1_in_6_valid,
  input        io_data_1_in_6_bits_valid,
  input  [7:0] io_data_1_in_6_bits_bits,
  input        io_data_1_in_7_valid,
  input        io_data_1_in_7_bits_valid,
  input  [7:0] io_data_1_in_7_bits_bits,
  input        io_data_1_in_8_valid,
  input        io_data_1_in_8_bits_valid,
  input  [7:0] io_data_1_in_8_bits_bits,
  input        io_data_1_in_9_valid,
  input        io_data_1_in_9_bits_valid,
  input  [7:0] io_data_1_in_9_bits_bits,
  input        io_data_1_in_10_valid,
  input        io_data_1_in_10_bits_valid,
  input  [7:0] io_data_1_in_10_bits_bits,
  input        io_data_1_in_11_valid,
  input        io_data_1_in_11_bits_valid,
  input  [7:0] io_data_1_in_11_bits_bits,
  input        io_data_1_in_12_valid,
  input        io_data_1_in_12_bits_valid,
  input  [7:0] io_data_1_in_12_bits_bits,
  input        io_data_1_in_13_valid,
  input        io_data_1_in_13_bits_valid,
  input  [7:0] io_data_1_in_13_bits_bits,
  input        io_data_1_in_14_valid,
  input        io_data_1_in_14_bits_valid,
  input  [7:0] io_data_1_in_14_bits_bits,
  input        io_data_1_in_15_valid,
  input        io_data_1_in_15_bits_valid,
  input  [7:0] io_data_1_in_15_bits_bits,
  output       io_data_0_out_0_valid,
  output [7:0] io_data_0_out_0_bits,
  output       io_data_0_out_1_valid,
  output [7:0] io_data_0_out_1_bits,
  output       io_data_0_out_2_valid,
  output [7:0] io_data_0_out_2_bits,
  output       io_data_0_out_3_valid,
  output [7:0] io_data_0_out_3_bits,
  output       io_data_0_out_4_valid,
  output [7:0] io_data_0_out_4_bits,
  output       io_data_0_out_5_valid,
  output [7:0] io_data_0_out_5_bits,
  output       io_data_0_out_6_valid,
  output [7:0] io_data_0_out_6_bits,
  output       io_data_0_out_7_valid,
  output [7:0] io_data_0_out_7_bits,
  output       io_data_0_out_8_valid,
  output [7:0] io_data_0_out_8_bits,
  output       io_data_0_out_9_valid,
  output [7:0] io_data_0_out_9_bits,
  output       io_data_0_out_10_valid,
  output [7:0] io_data_0_out_10_bits,
  output       io_data_0_out_11_valid,
  output [7:0] io_data_0_out_11_bits,
  output       io_data_0_out_12_valid,
  output [7:0] io_data_0_out_12_bits,
  output       io_data_0_out_13_valid,
  output [7:0] io_data_0_out_13_bits,
  output       io_data_0_out_14_valid,
  output [7:0] io_data_0_out_14_bits,
  output       io_data_0_out_15_valid,
  output [7:0] io_data_0_out_15_bits,
  input        io_exec_valid,
  input        io_out_valid
);
  wire  MultiDimTime_clock; // @[pearray.scala 63:25]
  wire  MultiDimTime_reset; // @[pearray.scala 63:25]
  wire  MultiDimTime_io_in; // @[pearray.scala 63:25]
  wire [1:0] MultiDimTime_io_out_0; // @[pearray.scala 63:25]
  wire [1:0] MultiDimTime_io_out_1; // @[pearray.scala 63:25]
  wire [17:0] MultiDimTime_io_index_0; // @[pearray.scala 63:25]
  wire [17:0] MultiDimTime_io_index_1; // @[pearray.scala 63:25]
  wire  PE_clock; // @[pearray.scala 101:13]
  wire  PE_reset; // @[pearray.scala 101:13]
  wire [7:0] PE_io_data_2_in_bits; // @[pearray.scala 101:13]
  wire [7:0] PE_io_data_2_out_bits; // @[pearray.scala 101:13]
  wire  PE_io_data_1_in_valid; // @[pearray.scala 101:13]
  wire [7:0] PE_io_data_1_in_bits; // @[pearray.scala 101:13]
  wire  PE_io_data_1_out_valid; // @[pearray.scala 101:13]
  wire [7:0] PE_io_data_1_out_bits; // @[pearray.scala 101:13]
  wire  PE_io_data_0_in_valid; // @[pearray.scala 101:13]
  wire [7:0] PE_io_data_0_in_bits; // @[pearray.scala 101:13]
  wire  PE_io_data_0_out_valid; // @[pearray.scala 101:13]
  wire [7:0] PE_io_data_0_out_bits; // @[pearray.scala 101:13]
  wire  PE_io_sig_stat2trans; // @[pearray.scala 101:13]
  wire  PE_1_clock; // @[pearray.scala 101:13]
  wire  PE_1_reset; // @[pearray.scala 101:13]
  wire [7:0] PE_1_io_data_2_in_bits; // @[pearray.scala 101:13]
  wire [7:0] PE_1_io_data_2_out_bits; // @[pearray.scala 101:13]
  wire  PE_1_io_data_1_in_valid; // @[pearray.scala 101:13]
  wire [7:0] PE_1_io_data_1_in_bits; // @[pearray.scala 101:13]
  wire  PE_1_io_data_1_out_valid; // @[pearray.scala 101:13]
  wire [7:0] PE_1_io_data_1_out_bits; // @[pearray.scala 101:13]
  wire  PE_1_io_data_0_in_valid; // @[pearray.scala 101:13]
  wire [7:0] PE_1_io_data_0_in_bits; // @[pearray.scala 101:13]
  wire  PE_1_io_data_0_out_valid; // @[pearray.scala 101:13]
  wire [7:0] PE_1_io_data_0_out_bits; // @[pearray.scala 101:13]
  wire  PE_1_io_sig_stat2trans; // @[pearray.scala 101:13]
  wire  PE_2_clock; // @[pearray.scala 101:13]
  wire  PE_2_reset; // @[pearray.scala 101:13]
  wire [7:0] PE_2_io_data_2_in_bits; // @[pearray.scala 101:13]
  wire [7:0] PE_2_io_data_2_out_bits; // @[pearray.scala 101:13]
  wire  PE_2_io_data_1_in_valid; // @[pearray.scala 101:13]
  wire [7:0] PE_2_io_data_1_in_bits; // @[pearray.scala 101:13]
  wire  PE_2_io_data_1_out_valid; // @[pearray.scala 101:13]
  wire [7:0] PE_2_io_data_1_out_bits; // @[pearray.scala 101:13]
  wire  PE_2_io_data_0_in_valid; // @[pearray.scala 101:13]
  wire [7:0] PE_2_io_data_0_in_bits; // @[pearray.scala 101:13]
  wire  PE_2_io_data_0_out_valid; // @[pearray.scala 101:13]
  wire [7:0] PE_2_io_data_0_out_bits; // @[pearray.scala 101:13]
  wire  PE_2_io_sig_stat2trans; // @[pearray.scala 101:13]
  wire  PE_3_clock; // @[pearray.scala 101:13]
  wire  PE_3_reset; // @[pearray.scala 101:13]
  wire [7:0] PE_3_io_data_2_in_bits; // @[pearray.scala 101:13]
  wire [7:0] PE_3_io_data_2_out_bits; // @[pearray.scala 101:13]
  wire  PE_3_io_data_1_in_valid; // @[pearray.scala 101:13]
  wire [7:0] PE_3_io_data_1_in_bits; // @[pearray.scala 101:13]
  wire  PE_3_io_data_1_out_valid; // @[pearray.scala 101:13]
  wire [7:0] PE_3_io_data_1_out_bits; // @[pearray.scala 101:13]
  wire  PE_3_io_data_0_in_valid; // @[pearray.scala 101:13]
  wire [7:0] PE_3_io_data_0_in_bits; // @[pearray.scala 101:13]
  wire  PE_3_io_data_0_out_valid; // @[pearray.scala 101:13]
  wire [7:0] PE_3_io_data_0_out_bits; // @[pearray.scala 101:13]
  wire  PE_3_io_sig_stat2trans; // @[pearray.scala 101:13]
  wire  PE_4_clock; // @[pearray.scala 101:13]
  wire  PE_4_reset; // @[pearray.scala 101:13]
  wire [7:0] PE_4_io_data_2_in_bits; // @[pearray.scala 101:13]
  wire [7:0] PE_4_io_data_2_out_bits; // @[pearray.scala 101:13]
  wire  PE_4_io_data_1_in_valid; // @[pearray.scala 101:13]
  wire [7:0] PE_4_io_data_1_in_bits; // @[pearray.scala 101:13]
  wire  PE_4_io_data_1_out_valid; // @[pearray.scala 101:13]
  wire [7:0] PE_4_io_data_1_out_bits; // @[pearray.scala 101:13]
  wire  PE_4_io_data_0_in_valid; // @[pearray.scala 101:13]
  wire [7:0] PE_4_io_data_0_in_bits; // @[pearray.scala 101:13]
  wire  PE_4_io_data_0_out_valid; // @[pearray.scala 101:13]
  wire [7:0] PE_4_io_data_0_out_bits; // @[pearray.scala 101:13]
  wire  PE_4_io_sig_stat2trans; // @[pearray.scala 101:13]
  wire  PE_5_clock; // @[pearray.scala 101:13]
  wire  PE_5_reset; // @[pearray.scala 101:13]
  wire [7:0] PE_5_io_data_2_in_bits; // @[pearray.scala 101:13]
  wire [7:0] PE_5_io_data_2_out_bits; // @[pearray.scala 101:13]
  wire  PE_5_io_data_1_in_valid; // @[pearray.scala 101:13]
  wire [7:0] PE_5_io_data_1_in_bits; // @[pearray.scala 101:13]
  wire  PE_5_io_data_1_out_valid; // @[pearray.scala 101:13]
  wire [7:0] PE_5_io_data_1_out_bits; // @[pearray.scala 101:13]
  wire  PE_5_io_data_0_in_valid; // @[pearray.scala 101:13]
  wire [7:0] PE_5_io_data_0_in_bits; // @[pearray.scala 101:13]
  wire  PE_5_io_data_0_out_valid; // @[pearray.scala 101:13]
  wire [7:0] PE_5_io_data_0_out_bits; // @[pearray.scala 101:13]
  wire  PE_5_io_sig_stat2trans; // @[pearray.scala 101:13]
  wire  PE_6_clock; // @[pearray.scala 101:13]
  wire  PE_6_reset; // @[pearray.scala 101:13]
  wire [7:0] PE_6_io_data_2_in_bits; // @[pearray.scala 101:13]
  wire [7:0] PE_6_io_data_2_out_bits; // @[pearray.scala 101:13]
  wire  PE_6_io_data_1_in_valid; // @[pearray.scala 101:13]
  wire [7:0] PE_6_io_data_1_in_bits; // @[pearray.scala 101:13]
  wire  PE_6_io_data_1_out_valid; // @[pearray.scala 101:13]
  wire [7:0] PE_6_io_data_1_out_bits; // @[pearray.scala 101:13]
  wire  PE_6_io_data_0_in_valid; // @[pearray.scala 101:13]
  wire [7:0] PE_6_io_data_0_in_bits; // @[pearray.scala 101:13]
  wire  PE_6_io_data_0_out_valid; // @[pearray.scala 101:13]
  wire [7:0] PE_6_io_data_0_out_bits; // @[pearray.scala 101:13]
  wire  PE_6_io_sig_stat2trans; // @[pearray.scala 101:13]
  wire  PE_7_clock; // @[pearray.scala 101:13]
  wire  PE_7_reset; // @[pearray.scala 101:13]
  wire [7:0] PE_7_io_data_2_in_bits; // @[pearray.scala 101:13]
  wire [7:0] PE_7_io_data_2_out_bits; // @[pearray.scala 101:13]
  wire  PE_7_io_data_1_in_valid; // @[pearray.scala 101:13]
  wire [7:0] PE_7_io_data_1_in_bits; // @[pearray.scala 101:13]
  wire  PE_7_io_data_1_out_valid; // @[pearray.scala 101:13]
  wire [7:0] PE_7_io_data_1_out_bits; // @[pearray.scala 101:13]
  wire  PE_7_io_data_0_in_valid; // @[pearray.scala 101:13]
  wire [7:0] PE_7_io_data_0_in_bits; // @[pearray.scala 101:13]
  wire  PE_7_io_data_0_out_valid; // @[pearray.scala 101:13]
  wire [7:0] PE_7_io_data_0_out_bits; // @[pearray.scala 101:13]
  wire  PE_7_io_sig_stat2trans; // @[pearray.scala 101:13]
  wire  PE_8_clock; // @[pearray.scala 101:13]
  wire  PE_8_reset; // @[pearray.scala 101:13]
  wire [7:0] PE_8_io_data_2_in_bits; // @[pearray.scala 101:13]
  wire [7:0] PE_8_io_data_2_out_bits; // @[pearray.scala 101:13]
  wire  PE_8_io_data_1_in_valid; // @[pearray.scala 101:13]
  wire [7:0] PE_8_io_data_1_in_bits; // @[pearray.scala 101:13]
  wire  PE_8_io_data_1_out_valid; // @[pearray.scala 101:13]
  wire [7:0] PE_8_io_data_1_out_bits; // @[pearray.scala 101:13]
  wire  PE_8_io_data_0_in_valid; // @[pearray.scala 101:13]
  wire [7:0] PE_8_io_data_0_in_bits; // @[pearray.scala 101:13]
  wire  PE_8_io_data_0_out_valid; // @[pearray.scala 101:13]
  wire [7:0] PE_8_io_data_0_out_bits; // @[pearray.scala 101:13]
  wire  PE_8_io_sig_stat2trans; // @[pearray.scala 101:13]
  wire  PE_9_clock; // @[pearray.scala 101:13]
  wire  PE_9_reset; // @[pearray.scala 101:13]
  wire [7:0] PE_9_io_data_2_in_bits; // @[pearray.scala 101:13]
  wire [7:0] PE_9_io_data_2_out_bits; // @[pearray.scala 101:13]
  wire  PE_9_io_data_1_in_valid; // @[pearray.scala 101:13]
  wire [7:0] PE_9_io_data_1_in_bits; // @[pearray.scala 101:13]
  wire  PE_9_io_data_1_out_valid; // @[pearray.scala 101:13]
  wire [7:0] PE_9_io_data_1_out_bits; // @[pearray.scala 101:13]
  wire  PE_9_io_data_0_in_valid; // @[pearray.scala 101:13]
  wire [7:0] PE_9_io_data_0_in_bits; // @[pearray.scala 101:13]
  wire  PE_9_io_data_0_out_valid; // @[pearray.scala 101:13]
  wire [7:0] PE_9_io_data_0_out_bits; // @[pearray.scala 101:13]
  wire  PE_9_io_sig_stat2trans; // @[pearray.scala 101:13]
  wire  PE_10_clock; // @[pearray.scala 101:13]
  wire  PE_10_reset; // @[pearray.scala 101:13]
  wire [7:0] PE_10_io_data_2_in_bits; // @[pearray.scala 101:13]
  wire [7:0] PE_10_io_data_2_out_bits; // @[pearray.scala 101:13]
  wire  PE_10_io_data_1_in_valid; // @[pearray.scala 101:13]
  wire [7:0] PE_10_io_data_1_in_bits; // @[pearray.scala 101:13]
  wire  PE_10_io_data_1_out_valid; // @[pearray.scala 101:13]
  wire [7:0] PE_10_io_data_1_out_bits; // @[pearray.scala 101:13]
  wire  PE_10_io_data_0_in_valid; // @[pearray.scala 101:13]
  wire [7:0] PE_10_io_data_0_in_bits; // @[pearray.scala 101:13]
  wire  PE_10_io_data_0_out_valid; // @[pearray.scala 101:13]
  wire [7:0] PE_10_io_data_0_out_bits; // @[pearray.scala 101:13]
  wire  PE_10_io_sig_stat2trans; // @[pearray.scala 101:13]
  wire  PE_11_clock; // @[pearray.scala 101:13]
  wire  PE_11_reset; // @[pearray.scala 101:13]
  wire [7:0] PE_11_io_data_2_in_bits; // @[pearray.scala 101:13]
  wire [7:0] PE_11_io_data_2_out_bits; // @[pearray.scala 101:13]
  wire  PE_11_io_data_1_in_valid; // @[pearray.scala 101:13]
  wire [7:0] PE_11_io_data_1_in_bits; // @[pearray.scala 101:13]
  wire  PE_11_io_data_1_out_valid; // @[pearray.scala 101:13]
  wire [7:0] PE_11_io_data_1_out_bits; // @[pearray.scala 101:13]
  wire  PE_11_io_data_0_in_valid; // @[pearray.scala 101:13]
  wire [7:0] PE_11_io_data_0_in_bits; // @[pearray.scala 101:13]
  wire  PE_11_io_data_0_out_valid; // @[pearray.scala 101:13]
  wire [7:0] PE_11_io_data_0_out_bits; // @[pearray.scala 101:13]
  wire  PE_11_io_sig_stat2trans; // @[pearray.scala 101:13]
  wire  PE_12_clock; // @[pearray.scala 101:13]
  wire  PE_12_reset; // @[pearray.scala 101:13]
  wire [7:0] PE_12_io_data_2_in_bits; // @[pearray.scala 101:13]
  wire [7:0] PE_12_io_data_2_out_bits; // @[pearray.scala 101:13]
  wire  PE_12_io_data_1_in_valid; // @[pearray.scala 101:13]
  wire [7:0] PE_12_io_data_1_in_bits; // @[pearray.scala 101:13]
  wire  PE_12_io_data_1_out_valid; // @[pearray.scala 101:13]
  wire [7:0] PE_12_io_data_1_out_bits; // @[pearray.scala 101:13]
  wire  PE_12_io_data_0_in_valid; // @[pearray.scala 101:13]
  wire [7:0] PE_12_io_data_0_in_bits; // @[pearray.scala 101:13]
  wire  PE_12_io_data_0_out_valid; // @[pearray.scala 101:13]
  wire [7:0] PE_12_io_data_0_out_bits; // @[pearray.scala 101:13]
  wire  PE_12_io_sig_stat2trans; // @[pearray.scala 101:13]
  wire  PE_13_clock; // @[pearray.scala 101:13]
  wire  PE_13_reset; // @[pearray.scala 101:13]
  wire [7:0] PE_13_io_data_2_in_bits; // @[pearray.scala 101:13]
  wire [7:0] PE_13_io_data_2_out_bits; // @[pearray.scala 101:13]
  wire  PE_13_io_data_1_in_valid; // @[pearray.scala 101:13]
  wire [7:0] PE_13_io_data_1_in_bits; // @[pearray.scala 101:13]
  wire  PE_13_io_data_1_out_valid; // @[pearray.scala 101:13]
  wire [7:0] PE_13_io_data_1_out_bits; // @[pearray.scala 101:13]
  wire  PE_13_io_data_0_in_valid; // @[pearray.scala 101:13]
  wire [7:0] PE_13_io_data_0_in_bits; // @[pearray.scala 101:13]
  wire  PE_13_io_data_0_out_valid; // @[pearray.scala 101:13]
  wire [7:0] PE_13_io_data_0_out_bits; // @[pearray.scala 101:13]
  wire  PE_13_io_sig_stat2trans; // @[pearray.scala 101:13]
  wire  PE_14_clock; // @[pearray.scala 101:13]
  wire  PE_14_reset; // @[pearray.scala 101:13]
  wire [7:0] PE_14_io_data_2_in_bits; // @[pearray.scala 101:13]
  wire [7:0] PE_14_io_data_2_out_bits; // @[pearray.scala 101:13]
  wire  PE_14_io_data_1_in_valid; // @[pearray.scala 101:13]
  wire [7:0] PE_14_io_data_1_in_bits; // @[pearray.scala 101:13]
  wire  PE_14_io_data_1_out_valid; // @[pearray.scala 101:13]
  wire [7:0] PE_14_io_data_1_out_bits; // @[pearray.scala 101:13]
  wire  PE_14_io_data_0_in_valid; // @[pearray.scala 101:13]
  wire [7:0] PE_14_io_data_0_in_bits; // @[pearray.scala 101:13]
  wire  PE_14_io_data_0_out_valid; // @[pearray.scala 101:13]
  wire [7:0] PE_14_io_data_0_out_bits; // @[pearray.scala 101:13]
  wire  PE_14_io_sig_stat2trans; // @[pearray.scala 101:13]
  wire  PE_15_clock; // @[pearray.scala 101:13]
  wire  PE_15_reset; // @[pearray.scala 101:13]
  wire [7:0] PE_15_io_data_2_in_bits; // @[pearray.scala 101:13]
  wire [7:0] PE_15_io_data_2_out_bits; // @[pearray.scala 101:13]
  wire  PE_15_io_data_1_in_valid; // @[pearray.scala 101:13]
  wire [7:0] PE_15_io_data_1_in_bits; // @[pearray.scala 101:13]
  wire  PE_15_io_data_1_out_valid; // @[pearray.scala 101:13]
  wire [7:0] PE_15_io_data_1_out_bits; // @[pearray.scala 101:13]
  wire  PE_15_io_data_0_in_valid; // @[pearray.scala 101:13]
  wire [7:0] PE_15_io_data_0_in_bits; // @[pearray.scala 101:13]
  wire  PE_15_io_data_0_out_valid; // @[pearray.scala 101:13]
  wire [7:0] PE_15_io_data_0_out_bits; // @[pearray.scala 101:13]
  wire  PE_15_io_sig_stat2trans; // @[pearray.scala 101:13]
  wire  PE_16_clock; // @[pearray.scala 101:13]
  wire  PE_16_reset; // @[pearray.scala 101:13]
  wire [7:0] PE_16_io_data_2_in_bits; // @[pearray.scala 101:13]
  wire [7:0] PE_16_io_data_2_out_bits; // @[pearray.scala 101:13]
  wire  PE_16_io_data_1_in_valid; // @[pearray.scala 101:13]
  wire [7:0] PE_16_io_data_1_in_bits; // @[pearray.scala 101:13]
  wire  PE_16_io_data_1_out_valid; // @[pearray.scala 101:13]
  wire [7:0] PE_16_io_data_1_out_bits; // @[pearray.scala 101:13]
  wire  PE_16_io_data_0_in_valid; // @[pearray.scala 101:13]
  wire [7:0] PE_16_io_data_0_in_bits; // @[pearray.scala 101:13]
  wire  PE_16_io_data_0_out_valid; // @[pearray.scala 101:13]
  wire [7:0] PE_16_io_data_0_out_bits; // @[pearray.scala 101:13]
  wire  PE_16_io_sig_stat2trans; // @[pearray.scala 101:13]
  wire  PE_17_clock; // @[pearray.scala 101:13]
  wire  PE_17_reset; // @[pearray.scala 101:13]
  wire [7:0] PE_17_io_data_2_in_bits; // @[pearray.scala 101:13]
  wire [7:0] PE_17_io_data_2_out_bits; // @[pearray.scala 101:13]
  wire  PE_17_io_data_1_in_valid; // @[pearray.scala 101:13]
  wire [7:0] PE_17_io_data_1_in_bits; // @[pearray.scala 101:13]
  wire  PE_17_io_data_1_out_valid; // @[pearray.scala 101:13]
  wire [7:0] PE_17_io_data_1_out_bits; // @[pearray.scala 101:13]
  wire  PE_17_io_data_0_in_valid; // @[pearray.scala 101:13]
  wire [7:0] PE_17_io_data_0_in_bits; // @[pearray.scala 101:13]
  wire  PE_17_io_data_0_out_valid; // @[pearray.scala 101:13]
  wire [7:0] PE_17_io_data_0_out_bits; // @[pearray.scala 101:13]
  wire  PE_17_io_sig_stat2trans; // @[pearray.scala 101:13]
  wire  PE_18_clock; // @[pearray.scala 101:13]
  wire  PE_18_reset; // @[pearray.scala 101:13]
  wire [7:0] PE_18_io_data_2_in_bits; // @[pearray.scala 101:13]
  wire [7:0] PE_18_io_data_2_out_bits; // @[pearray.scala 101:13]
  wire  PE_18_io_data_1_in_valid; // @[pearray.scala 101:13]
  wire [7:0] PE_18_io_data_1_in_bits; // @[pearray.scala 101:13]
  wire  PE_18_io_data_1_out_valid; // @[pearray.scala 101:13]
  wire [7:0] PE_18_io_data_1_out_bits; // @[pearray.scala 101:13]
  wire  PE_18_io_data_0_in_valid; // @[pearray.scala 101:13]
  wire [7:0] PE_18_io_data_0_in_bits; // @[pearray.scala 101:13]
  wire  PE_18_io_data_0_out_valid; // @[pearray.scala 101:13]
  wire [7:0] PE_18_io_data_0_out_bits; // @[pearray.scala 101:13]
  wire  PE_18_io_sig_stat2trans; // @[pearray.scala 101:13]
  wire  PE_19_clock; // @[pearray.scala 101:13]
  wire  PE_19_reset; // @[pearray.scala 101:13]
  wire [7:0] PE_19_io_data_2_in_bits; // @[pearray.scala 101:13]
  wire [7:0] PE_19_io_data_2_out_bits; // @[pearray.scala 101:13]
  wire  PE_19_io_data_1_in_valid; // @[pearray.scala 101:13]
  wire [7:0] PE_19_io_data_1_in_bits; // @[pearray.scala 101:13]
  wire  PE_19_io_data_1_out_valid; // @[pearray.scala 101:13]
  wire [7:0] PE_19_io_data_1_out_bits; // @[pearray.scala 101:13]
  wire  PE_19_io_data_0_in_valid; // @[pearray.scala 101:13]
  wire [7:0] PE_19_io_data_0_in_bits; // @[pearray.scala 101:13]
  wire  PE_19_io_data_0_out_valid; // @[pearray.scala 101:13]
  wire [7:0] PE_19_io_data_0_out_bits; // @[pearray.scala 101:13]
  wire  PE_19_io_sig_stat2trans; // @[pearray.scala 101:13]
  wire  PE_20_clock; // @[pearray.scala 101:13]
  wire  PE_20_reset; // @[pearray.scala 101:13]
  wire [7:0] PE_20_io_data_2_in_bits; // @[pearray.scala 101:13]
  wire [7:0] PE_20_io_data_2_out_bits; // @[pearray.scala 101:13]
  wire  PE_20_io_data_1_in_valid; // @[pearray.scala 101:13]
  wire [7:0] PE_20_io_data_1_in_bits; // @[pearray.scala 101:13]
  wire  PE_20_io_data_1_out_valid; // @[pearray.scala 101:13]
  wire [7:0] PE_20_io_data_1_out_bits; // @[pearray.scala 101:13]
  wire  PE_20_io_data_0_in_valid; // @[pearray.scala 101:13]
  wire [7:0] PE_20_io_data_0_in_bits; // @[pearray.scala 101:13]
  wire  PE_20_io_data_0_out_valid; // @[pearray.scala 101:13]
  wire [7:0] PE_20_io_data_0_out_bits; // @[pearray.scala 101:13]
  wire  PE_20_io_sig_stat2trans; // @[pearray.scala 101:13]
  wire  PE_21_clock; // @[pearray.scala 101:13]
  wire  PE_21_reset; // @[pearray.scala 101:13]
  wire [7:0] PE_21_io_data_2_in_bits; // @[pearray.scala 101:13]
  wire [7:0] PE_21_io_data_2_out_bits; // @[pearray.scala 101:13]
  wire  PE_21_io_data_1_in_valid; // @[pearray.scala 101:13]
  wire [7:0] PE_21_io_data_1_in_bits; // @[pearray.scala 101:13]
  wire  PE_21_io_data_1_out_valid; // @[pearray.scala 101:13]
  wire [7:0] PE_21_io_data_1_out_bits; // @[pearray.scala 101:13]
  wire  PE_21_io_data_0_in_valid; // @[pearray.scala 101:13]
  wire [7:0] PE_21_io_data_0_in_bits; // @[pearray.scala 101:13]
  wire  PE_21_io_data_0_out_valid; // @[pearray.scala 101:13]
  wire [7:0] PE_21_io_data_0_out_bits; // @[pearray.scala 101:13]
  wire  PE_21_io_sig_stat2trans; // @[pearray.scala 101:13]
  wire  PE_22_clock; // @[pearray.scala 101:13]
  wire  PE_22_reset; // @[pearray.scala 101:13]
  wire [7:0] PE_22_io_data_2_in_bits; // @[pearray.scala 101:13]
  wire [7:0] PE_22_io_data_2_out_bits; // @[pearray.scala 101:13]
  wire  PE_22_io_data_1_in_valid; // @[pearray.scala 101:13]
  wire [7:0] PE_22_io_data_1_in_bits; // @[pearray.scala 101:13]
  wire  PE_22_io_data_1_out_valid; // @[pearray.scala 101:13]
  wire [7:0] PE_22_io_data_1_out_bits; // @[pearray.scala 101:13]
  wire  PE_22_io_data_0_in_valid; // @[pearray.scala 101:13]
  wire [7:0] PE_22_io_data_0_in_bits; // @[pearray.scala 101:13]
  wire  PE_22_io_data_0_out_valid; // @[pearray.scala 101:13]
  wire [7:0] PE_22_io_data_0_out_bits; // @[pearray.scala 101:13]
  wire  PE_22_io_sig_stat2trans; // @[pearray.scala 101:13]
  wire  PE_23_clock; // @[pearray.scala 101:13]
  wire  PE_23_reset; // @[pearray.scala 101:13]
  wire [7:0] PE_23_io_data_2_in_bits; // @[pearray.scala 101:13]
  wire [7:0] PE_23_io_data_2_out_bits; // @[pearray.scala 101:13]
  wire  PE_23_io_data_1_in_valid; // @[pearray.scala 101:13]
  wire [7:0] PE_23_io_data_1_in_bits; // @[pearray.scala 101:13]
  wire  PE_23_io_data_1_out_valid; // @[pearray.scala 101:13]
  wire [7:0] PE_23_io_data_1_out_bits; // @[pearray.scala 101:13]
  wire  PE_23_io_data_0_in_valid; // @[pearray.scala 101:13]
  wire [7:0] PE_23_io_data_0_in_bits; // @[pearray.scala 101:13]
  wire  PE_23_io_data_0_out_valid; // @[pearray.scala 101:13]
  wire [7:0] PE_23_io_data_0_out_bits; // @[pearray.scala 101:13]
  wire  PE_23_io_sig_stat2trans; // @[pearray.scala 101:13]
  wire  PE_24_clock; // @[pearray.scala 101:13]
  wire  PE_24_reset; // @[pearray.scala 101:13]
  wire [7:0] PE_24_io_data_2_in_bits; // @[pearray.scala 101:13]
  wire [7:0] PE_24_io_data_2_out_bits; // @[pearray.scala 101:13]
  wire  PE_24_io_data_1_in_valid; // @[pearray.scala 101:13]
  wire [7:0] PE_24_io_data_1_in_bits; // @[pearray.scala 101:13]
  wire  PE_24_io_data_1_out_valid; // @[pearray.scala 101:13]
  wire [7:0] PE_24_io_data_1_out_bits; // @[pearray.scala 101:13]
  wire  PE_24_io_data_0_in_valid; // @[pearray.scala 101:13]
  wire [7:0] PE_24_io_data_0_in_bits; // @[pearray.scala 101:13]
  wire  PE_24_io_data_0_out_valid; // @[pearray.scala 101:13]
  wire [7:0] PE_24_io_data_0_out_bits; // @[pearray.scala 101:13]
  wire  PE_24_io_sig_stat2trans; // @[pearray.scala 101:13]
  wire  PE_25_clock; // @[pearray.scala 101:13]
  wire  PE_25_reset; // @[pearray.scala 101:13]
  wire [7:0] PE_25_io_data_2_in_bits; // @[pearray.scala 101:13]
  wire [7:0] PE_25_io_data_2_out_bits; // @[pearray.scala 101:13]
  wire  PE_25_io_data_1_in_valid; // @[pearray.scala 101:13]
  wire [7:0] PE_25_io_data_1_in_bits; // @[pearray.scala 101:13]
  wire  PE_25_io_data_1_out_valid; // @[pearray.scala 101:13]
  wire [7:0] PE_25_io_data_1_out_bits; // @[pearray.scala 101:13]
  wire  PE_25_io_data_0_in_valid; // @[pearray.scala 101:13]
  wire [7:0] PE_25_io_data_0_in_bits; // @[pearray.scala 101:13]
  wire  PE_25_io_data_0_out_valid; // @[pearray.scala 101:13]
  wire [7:0] PE_25_io_data_0_out_bits; // @[pearray.scala 101:13]
  wire  PE_25_io_sig_stat2trans; // @[pearray.scala 101:13]
  wire  PE_26_clock; // @[pearray.scala 101:13]
  wire  PE_26_reset; // @[pearray.scala 101:13]
  wire [7:0] PE_26_io_data_2_in_bits; // @[pearray.scala 101:13]
  wire [7:0] PE_26_io_data_2_out_bits; // @[pearray.scala 101:13]
  wire  PE_26_io_data_1_in_valid; // @[pearray.scala 101:13]
  wire [7:0] PE_26_io_data_1_in_bits; // @[pearray.scala 101:13]
  wire  PE_26_io_data_1_out_valid; // @[pearray.scala 101:13]
  wire [7:0] PE_26_io_data_1_out_bits; // @[pearray.scala 101:13]
  wire  PE_26_io_data_0_in_valid; // @[pearray.scala 101:13]
  wire [7:0] PE_26_io_data_0_in_bits; // @[pearray.scala 101:13]
  wire  PE_26_io_data_0_out_valid; // @[pearray.scala 101:13]
  wire [7:0] PE_26_io_data_0_out_bits; // @[pearray.scala 101:13]
  wire  PE_26_io_sig_stat2trans; // @[pearray.scala 101:13]
  wire  PE_27_clock; // @[pearray.scala 101:13]
  wire  PE_27_reset; // @[pearray.scala 101:13]
  wire [7:0] PE_27_io_data_2_in_bits; // @[pearray.scala 101:13]
  wire [7:0] PE_27_io_data_2_out_bits; // @[pearray.scala 101:13]
  wire  PE_27_io_data_1_in_valid; // @[pearray.scala 101:13]
  wire [7:0] PE_27_io_data_1_in_bits; // @[pearray.scala 101:13]
  wire  PE_27_io_data_1_out_valid; // @[pearray.scala 101:13]
  wire [7:0] PE_27_io_data_1_out_bits; // @[pearray.scala 101:13]
  wire  PE_27_io_data_0_in_valid; // @[pearray.scala 101:13]
  wire [7:0] PE_27_io_data_0_in_bits; // @[pearray.scala 101:13]
  wire  PE_27_io_data_0_out_valid; // @[pearray.scala 101:13]
  wire [7:0] PE_27_io_data_0_out_bits; // @[pearray.scala 101:13]
  wire  PE_27_io_sig_stat2trans; // @[pearray.scala 101:13]
  wire  PE_28_clock; // @[pearray.scala 101:13]
  wire  PE_28_reset; // @[pearray.scala 101:13]
  wire [7:0] PE_28_io_data_2_in_bits; // @[pearray.scala 101:13]
  wire [7:0] PE_28_io_data_2_out_bits; // @[pearray.scala 101:13]
  wire  PE_28_io_data_1_in_valid; // @[pearray.scala 101:13]
  wire [7:0] PE_28_io_data_1_in_bits; // @[pearray.scala 101:13]
  wire  PE_28_io_data_1_out_valid; // @[pearray.scala 101:13]
  wire [7:0] PE_28_io_data_1_out_bits; // @[pearray.scala 101:13]
  wire  PE_28_io_data_0_in_valid; // @[pearray.scala 101:13]
  wire [7:0] PE_28_io_data_0_in_bits; // @[pearray.scala 101:13]
  wire  PE_28_io_data_0_out_valid; // @[pearray.scala 101:13]
  wire [7:0] PE_28_io_data_0_out_bits; // @[pearray.scala 101:13]
  wire  PE_28_io_sig_stat2trans; // @[pearray.scala 101:13]
  wire  PE_29_clock; // @[pearray.scala 101:13]
  wire  PE_29_reset; // @[pearray.scala 101:13]
  wire [7:0] PE_29_io_data_2_in_bits; // @[pearray.scala 101:13]
  wire [7:0] PE_29_io_data_2_out_bits; // @[pearray.scala 101:13]
  wire  PE_29_io_data_1_in_valid; // @[pearray.scala 101:13]
  wire [7:0] PE_29_io_data_1_in_bits; // @[pearray.scala 101:13]
  wire  PE_29_io_data_1_out_valid; // @[pearray.scala 101:13]
  wire [7:0] PE_29_io_data_1_out_bits; // @[pearray.scala 101:13]
  wire  PE_29_io_data_0_in_valid; // @[pearray.scala 101:13]
  wire [7:0] PE_29_io_data_0_in_bits; // @[pearray.scala 101:13]
  wire  PE_29_io_data_0_out_valid; // @[pearray.scala 101:13]
  wire [7:0] PE_29_io_data_0_out_bits; // @[pearray.scala 101:13]
  wire  PE_29_io_sig_stat2trans; // @[pearray.scala 101:13]
  wire  PE_30_clock; // @[pearray.scala 101:13]
  wire  PE_30_reset; // @[pearray.scala 101:13]
  wire [7:0] PE_30_io_data_2_in_bits; // @[pearray.scala 101:13]
  wire [7:0] PE_30_io_data_2_out_bits; // @[pearray.scala 101:13]
  wire  PE_30_io_data_1_in_valid; // @[pearray.scala 101:13]
  wire [7:0] PE_30_io_data_1_in_bits; // @[pearray.scala 101:13]
  wire  PE_30_io_data_1_out_valid; // @[pearray.scala 101:13]
  wire [7:0] PE_30_io_data_1_out_bits; // @[pearray.scala 101:13]
  wire  PE_30_io_data_0_in_valid; // @[pearray.scala 101:13]
  wire [7:0] PE_30_io_data_0_in_bits; // @[pearray.scala 101:13]
  wire  PE_30_io_data_0_out_valid; // @[pearray.scala 101:13]
  wire [7:0] PE_30_io_data_0_out_bits; // @[pearray.scala 101:13]
  wire  PE_30_io_sig_stat2trans; // @[pearray.scala 101:13]
  wire  PE_31_clock; // @[pearray.scala 101:13]
  wire  PE_31_reset; // @[pearray.scala 101:13]
  wire [7:0] PE_31_io_data_2_in_bits; // @[pearray.scala 101:13]
  wire [7:0] PE_31_io_data_2_out_bits; // @[pearray.scala 101:13]
  wire  PE_31_io_data_1_in_valid; // @[pearray.scala 101:13]
  wire [7:0] PE_31_io_data_1_in_bits; // @[pearray.scala 101:13]
  wire  PE_31_io_data_1_out_valid; // @[pearray.scala 101:13]
  wire [7:0] PE_31_io_data_1_out_bits; // @[pearray.scala 101:13]
  wire  PE_31_io_data_0_in_valid; // @[pearray.scala 101:13]
  wire [7:0] PE_31_io_data_0_in_bits; // @[pearray.scala 101:13]
  wire  PE_31_io_data_0_out_valid; // @[pearray.scala 101:13]
  wire [7:0] PE_31_io_data_0_out_bits; // @[pearray.scala 101:13]
  wire  PE_31_io_sig_stat2trans; // @[pearray.scala 101:13]
  wire  PE_32_clock; // @[pearray.scala 101:13]
  wire  PE_32_reset; // @[pearray.scala 101:13]
  wire [7:0] PE_32_io_data_2_in_bits; // @[pearray.scala 101:13]
  wire [7:0] PE_32_io_data_2_out_bits; // @[pearray.scala 101:13]
  wire  PE_32_io_data_1_in_valid; // @[pearray.scala 101:13]
  wire [7:0] PE_32_io_data_1_in_bits; // @[pearray.scala 101:13]
  wire  PE_32_io_data_1_out_valid; // @[pearray.scala 101:13]
  wire [7:0] PE_32_io_data_1_out_bits; // @[pearray.scala 101:13]
  wire  PE_32_io_data_0_in_valid; // @[pearray.scala 101:13]
  wire [7:0] PE_32_io_data_0_in_bits; // @[pearray.scala 101:13]
  wire  PE_32_io_data_0_out_valid; // @[pearray.scala 101:13]
  wire [7:0] PE_32_io_data_0_out_bits; // @[pearray.scala 101:13]
  wire  PE_32_io_sig_stat2trans; // @[pearray.scala 101:13]
  wire  PE_33_clock; // @[pearray.scala 101:13]
  wire  PE_33_reset; // @[pearray.scala 101:13]
  wire [7:0] PE_33_io_data_2_in_bits; // @[pearray.scala 101:13]
  wire [7:0] PE_33_io_data_2_out_bits; // @[pearray.scala 101:13]
  wire  PE_33_io_data_1_in_valid; // @[pearray.scala 101:13]
  wire [7:0] PE_33_io_data_1_in_bits; // @[pearray.scala 101:13]
  wire  PE_33_io_data_1_out_valid; // @[pearray.scala 101:13]
  wire [7:0] PE_33_io_data_1_out_bits; // @[pearray.scala 101:13]
  wire  PE_33_io_data_0_in_valid; // @[pearray.scala 101:13]
  wire [7:0] PE_33_io_data_0_in_bits; // @[pearray.scala 101:13]
  wire  PE_33_io_data_0_out_valid; // @[pearray.scala 101:13]
  wire [7:0] PE_33_io_data_0_out_bits; // @[pearray.scala 101:13]
  wire  PE_33_io_sig_stat2trans; // @[pearray.scala 101:13]
  wire  PE_34_clock; // @[pearray.scala 101:13]
  wire  PE_34_reset; // @[pearray.scala 101:13]
  wire [7:0] PE_34_io_data_2_in_bits; // @[pearray.scala 101:13]
  wire [7:0] PE_34_io_data_2_out_bits; // @[pearray.scala 101:13]
  wire  PE_34_io_data_1_in_valid; // @[pearray.scala 101:13]
  wire [7:0] PE_34_io_data_1_in_bits; // @[pearray.scala 101:13]
  wire  PE_34_io_data_1_out_valid; // @[pearray.scala 101:13]
  wire [7:0] PE_34_io_data_1_out_bits; // @[pearray.scala 101:13]
  wire  PE_34_io_data_0_in_valid; // @[pearray.scala 101:13]
  wire [7:0] PE_34_io_data_0_in_bits; // @[pearray.scala 101:13]
  wire  PE_34_io_data_0_out_valid; // @[pearray.scala 101:13]
  wire [7:0] PE_34_io_data_0_out_bits; // @[pearray.scala 101:13]
  wire  PE_34_io_sig_stat2trans; // @[pearray.scala 101:13]
  wire  PE_35_clock; // @[pearray.scala 101:13]
  wire  PE_35_reset; // @[pearray.scala 101:13]
  wire [7:0] PE_35_io_data_2_in_bits; // @[pearray.scala 101:13]
  wire [7:0] PE_35_io_data_2_out_bits; // @[pearray.scala 101:13]
  wire  PE_35_io_data_1_in_valid; // @[pearray.scala 101:13]
  wire [7:0] PE_35_io_data_1_in_bits; // @[pearray.scala 101:13]
  wire  PE_35_io_data_1_out_valid; // @[pearray.scala 101:13]
  wire [7:0] PE_35_io_data_1_out_bits; // @[pearray.scala 101:13]
  wire  PE_35_io_data_0_in_valid; // @[pearray.scala 101:13]
  wire [7:0] PE_35_io_data_0_in_bits; // @[pearray.scala 101:13]
  wire  PE_35_io_data_0_out_valid; // @[pearray.scala 101:13]
  wire [7:0] PE_35_io_data_0_out_bits; // @[pearray.scala 101:13]
  wire  PE_35_io_sig_stat2trans; // @[pearray.scala 101:13]
  wire  PE_36_clock; // @[pearray.scala 101:13]
  wire  PE_36_reset; // @[pearray.scala 101:13]
  wire [7:0] PE_36_io_data_2_in_bits; // @[pearray.scala 101:13]
  wire [7:0] PE_36_io_data_2_out_bits; // @[pearray.scala 101:13]
  wire  PE_36_io_data_1_in_valid; // @[pearray.scala 101:13]
  wire [7:0] PE_36_io_data_1_in_bits; // @[pearray.scala 101:13]
  wire  PE_36_io_data_1_out_valid; // @[pearray.scala 101:13]
  wire [7:0] PE_36_io_data_1_out_bits; // @[pearray.scala 101:13]
  wire  PE_36_io_data_0_in_valid; // @[pearray.scala 101:13]
  wire [7:0] PE_36_io_data_0_in_bits; // @[pearray.scala 101:13]
  wire  PE_36_io_data_0_out_valid; // @[pearray.scala 101:13]
  wire [7:0] PE_36_io_data_0_out_bits; // @[pearray.scala 101:13]
  wire  PE_36_io_sig_stat2trans; // @[pearray.scala 101:13]
  wire  PE_37_clock; // @[pearray.scala 101:13]
  wire  PE_37_reset; // @[pearray.scala 101:13]
  wire [7:0] PE_37_io_data_2_in_bits; // @[pearray.scala 101:13]
  wire [7:0] PE_37_io_data_2_out_bits; // @[pearray.scala 101:13]
  wire  PE_37_io_data_1_in_valid; // @[pearray.scala 101:13]
  wire [7:0] PE_37_io_data_1_in_bits; // @[pearray.scala 101:13]
  wire  PE_37_io_data_1_out_valid; // @[pearray.scala 101:13]
  wire [7:0] PE_37_io_data_1_out_bits; // @[pearray.scala 101:13]
  wire  PE_37_io_data_0_in_valid; // @[pearray.scala 101:13]
  wire [7:0] PE_37_io_data_0_in_bits; // @[pearray.scala 101:13]
  wire  PE_37_io_data_0_out_valid; // @[pearray.scala 101:13]
  wire [7:0] PE_37_io_data_0_out_bits; // @[pearray.scala 101:13]
  wire  PE_37_io_sig_stat2trans; // @[pearray.scala 101:13]
  wire  PE_38_clock; // @[pearray.scala 101:13]
  wire  PE_38_reset; // @[pearray.scala 101:13]
  wire [7:0] PE_38_io_data_2_in_bits; // @[pearray.scala 101:13]
  wire [7:0] PE_38_io_data_2_out_bits; // @[pearray.scala 101:13]
  wire  PE_38_io_data_1_in_valid; // @[pearray.scala 101:13]
  wire [7:0] PE_38_io_data_1_in_bits; // @[pearray.scala 101:13]
  wire  PE_38_io_data_1_out_valid; // @[pearray.scala 101:13]
  wire [7:0] PE_38_io_data_1_out_bits; // @[pearray.scala 101:13]
  wire  PE_38_io_data_0_in_valid; // @[pearray.scala 101:13]
  wire [7:0] PE_38_io_data_0_in_bits; // @[pearray.scala 101:13]
  wire  PE_38_io_data_0_out_valid; // @[pearray.scala 101:13]
  wire [7:0] PE_38_io_data_0_out_bits; // @[pearray.scala 101:13]
  wire  PE_38_io_sig_stat2trans; // @[pearray.scala 101:13]
  wire  PE_39_clock; // @[pearray.scala 101:13]
  wire  PE_39_reset; // @[pearray.scala 101:13]
  wire [7:0] PE_39_io_data_2_in_bits; // @[pearray.scala 101:13]
  wire [7:0] PE_39_io_data_2_out_bits; // @[pearray.scala 101:13]
  wire  PE_39_io_data_1_in_valid; // @[pearray.scala 101:13]
  wire [7:0] PE_39_io_data_1_in_bits; // @[pearray.scala 101:13]
  wire  PE_39_io_data_1_out_valid; // @[pearray.scala 101:13]
  wire [7:0] PE_39_io_data_1_out_bits; // @[pearray.scala 101:13]
  wire  PE_39_io_data_0_in_valid; // @[pearray.scala 101:13]
  wire [7:0] PE_39_io_data_0_in_bits; // @[pearray.scala 101:13]
  wire  PE_39_io_data_0_out_valid; // @[pearray.scala 101:13]
  wire [7:0] PE_39_io_data_0_out_bits; // @[pearray.scala 101:13]
  wire  PE_39_io_sig_stat2trans; // @[pearray.scala 101:13]
  wire  PE_40_clock; // @[pearray.scala 101:13]
  wire  PE_40_reset; // @[pearray.scala 101:13]
  wire [7:0] PE_40_io_data_2_in_bits; // @[pearray.scala 101:13]
  wire [7:0] PE_40_io_data_2_out_bits; // @[pearray.scala 101:13]
  wire  PE_40_io_data_1_in_valid; // @[pearray.scala 101:13]
  wire [7:0] PE_40_io_data_1_in_bits; // @[pearray.scala 101:13]
  wire  PE_40_io_data_1_out_valid; // @[pearray.scala 101:13]
  wire [7:0] PE_40_io_data_1_out_bits; // @[pearray.scala 101:13]
  wire  PE_40_io_data_0_in_valid; // @[pearray.scala 101:13]
  wire [7:0] PE_40_io_data_0_in_bits; // @[pearray.scala 101:13]
  wire  PE_40_io_data_0_out_valid; // @[pearray.scala 101:13]
  wire [7:0] PE_40_io_data_0_out_bits; // @[pearray.scala 101:13]
  wire  PE_40_io_sig_stat2trans; // @[pearray.scala 101:13]
  wire  PE_41_clock; // @[pearray.scala 101:13]
  wire  PE_41_reset; // @[pearray.scala 101:13]
  wire [7:0] PE_41_io_data_2_in_bits; // @[pearray.scala 101:13]
  wire [7:0] PE_41_io_data_2_out_bits; // @[pearray.scala 101:13]
  wire  PE_41_io_data_1_in_valid; // @[pearray.scala 101:13]
  wire [7:0] PE_41_io_data_1_in_bits; // @[pearray.scala 101:13]
  wire  PE_41_io_data_1_out_valid; // @[pearray.scala 101:13]
  wire [7:0] PE_41_io_data_1_out_bits; // @[pearray.scala 101:13]
  wire  PE_41_io_data_0_in_valid; // @[pearray.scala 101:13]
  wire [7:0] PE_41_io_data_0_in_bits; // @[pearray.scala 101:13]
  wire  PE_41_io_data_0_out_valid; // @[pearray.scala 101:13]
  wire [7:0] PE_41_io_data_0_out_bits; // @[pearray.scala 101:13]
  wire  PE_41_io_sig_stat2trans; // @[pearray.scala 101:13]
  wire  PE_42_clock; // @[pearray.scala 101:13]
  wire  PE_42_reset; // @[pearray.scala 101:13]
  wire [7:0] PE_42_io_data_2_in_bits; // @[pearray.scala 101:13]
  wire [7:0] PE_42_io_data_2_out_bits; // @[pearray.scala 101:13]
  wire  PE_42_io_data_1_in_valid; // @[pearray.scala 101:13]
  wire [7:0] PE_42_io_data_1_in_bits; // @[pearray.scala 101:13]
  wire  PE_42_io_data_1_out_valid; // @[pearray.scala 101:13]
  wire [7:0] PE_42_io_data_1_out_bits; // @[pearray.scala 101:13]
  wire  PE_42_io_data_0_in_valid; // @[pearray.scala 101:13]
  wire [7:0] PE_42_io_data_0_in_bits; // @[pearray.scala 101:13]
  wire  PE_42_io_data_0_out_valid; // @[pearray.scala 101:13]
  wire [7:0] PE_42_io_data_0_out_bits; // @[pearray.scala 101:13]
  wire  PE_42_io_sig_stat2trans; // @[pearray.scala 101:13]
  wire  PE_43_clock; // @[pearray.scala 101:13]
  wire  PE_43_reset; // @[pearray.scala 101:13]
  wire [7:0] PE_43_io_data_2_in_bits; // @[pearray.scala 101:13]
  wire [7:0] PE_43_io_data_2_out_bits; // @[pearray.scala 101:13]
  wire  PE_43_io_data_1_in_valid; // @[pearray.scala 101:13]
  wire [7:0] PE_43_io_data_1_in_bits; // @[pearray.scala 101:13]
  wire  PE_43_io_data_1_out_valid; // @[pearray.scala 101:13]
  wire [7:0] PE_43_io_data_1_out_bits; // @[pearray.scala 101:13]
  wire  PE_43_io_data_0_in_valid; // @[pearray.scala 101:13]
  wire [7:0] PE_43_io_data_0_in_bits; // @[pearray.scala 101:13]
  wire  PE_43_io_data_0_out_valid; // @[pearray.scala 101:13]
  wire [7:0] PE_43_io_data_0_out_bits; // @[pearray.scala 101:13]
  wire  PE_43_io_sig_stat2trans; // @[pearray.scala 101:13]
  wire  PE_44_clock; // @[pearray.scala 101:13]
  wire  PE_44_reset; // @[pearray.scala 101:13]
  wire [7:0] PE_44_io_data_2_in_bits; // @[pearray.scala 101:13]
  wire [7:0] PE_44_io_data_2_out_bits; // @[pearray.scala 101:13]
  wire  PE_44_io_data_1_in_valid; // @[pearray.scala 101:13]
  wire [7:0] PE_44_io_data_1_in_bits; // @[pearray.scala 101:13]
  wire  PE_44_io_data_1_out_valid; // @[pearray.scala 101:13]
  wire [7:0] PE_44_io_data_1_out_bits; // @[pearray.scala 101:13]
  wire  PE_44_io_data_0_in_valid; // @[pearray.scala 101:13]
  wire [7:0] PE_44_io_data_0_in_bits; // @[pearray.scala 101:13]
  wire  PE_44_io_data_0_out_valid; // @[pearray.scala 101:13]
  wire [7:0] PE_44_io_data_0_out_bits; // @[pearray.scala 101:13]
  wire  PE_44_io_sig_stat2trans; // @[pearray.scala 101:13]
  wire  PE_45_clock; // @[pearray.scala 101:13]
  wire  PE_45_reset; // @[pearray.scala 101:13]
  wire [7:0] PE_45_io_data_2_in_bits; // @[pearray.scala 101:13]
  wire [7:0] PE_45_io_data_2_out_bits; // @[pearray.scala 101:13]
  wire  PE_45_io_data_1_in_valid; // @[pearray.scala 101:13]
  wire [7:0] PE_45_io_data_1_in_bits; // @[pearray.scala 101:13]
  wire  PE_45_io_data_1_out_valid; // @[pearray.scala 101:13]
  wire [7:0] PE_45_io_data_1_out_bits; // @[pearray.scala 101:13]
  wire  PE_45_io_data_0_in_valid; // @[pearray.scala 101:13]
  wire [7:0] PE_45_io_data_0_in_bits; // @[pearray.scala 101:13]
  wire  PE_45_io_data_0_out_valid; // @[pearray.scala 101:13]
  wire [7:0] PE_45_io_data_0_out_bits; // @[pearray.scala 101:13]
  wire  PE_45_io_sig_stat2trans; // @[pearray.scala 101:13]
  wire  PE_46_clock; // @[pearray.scala 101:13]
  wire  PE_46_reset; // @[pearray.scala 101:13]
  wire [7:0] PE_46_io_data_2_in_bits; // @[pearray.scala 101:13]
  wire [7:0] PE_46_io_data_2_out_bits; // @[pearray.scala 101:13]
  wire  PE_46_io_data_1_in_valid; // @[pearray.scala 101:13]
  wire [7:0] PE_46_io_data_1_in_bits; // @[pearray.scala 101:13]
  wire  PE_46_io_data_1_out_valid; // @[pearray.scala 101:13]
  wire [7:0] PE_46_io_data_1_out_bits; // @[pearray.scala 101:13]
  wire  PE_46_io_data_0_in_valid; // @[pearray.scala 101:13]
  wire [7:0] PE_46_io_data_0_in_bits; // @[pearray.scala 101:13]
  wire  PE_46_io_data_0_out_valid; // @[pearray.scala 101:13]
  wire [7:0] PE_46_io_data_0_out_bits; // @[pearray.scala 101:13]
  wire  PE_46_io_sig_stat2trans; // @[pearray.scala 101:13]
  wire  PE_47_clock; // @[pearray.scala 101:13]
  wire  PE_47_reset; // @[pearray.scala 101:13]
  wire [7:0] PE_47_io_data_2_in_bits; // @[pearray.scala 101:13]
  wire [7:0] PE_47_io_data_2_out_bits; // @[pearray.scala 101:13]
  wire  PE_47_io_data_1_in_valid; // @[pearray.scala 101:13]
  wire [7:0] PE_47_io_data_1_in_bits; // @[pearray.scala 101:13]
  wire  PE_47_io_data_1_out_valid; // @[pearray.scala 101:13]
  wire [7:0] PE_47_io_data_1_out_bits; // @[pearray.scala 101:13]
  wire  PE_47_io_data_0_in_valid; // @[pearray.scala 101:13]
  wire [7:0] PE_47_io_data_0_in_bits; // @[pearray.scala 101:13]
  wire  PE_47_io_data_0_out_valid; // @[pearray.scala 101:13]
  wire [7:0] PE_47_io_data_0_out_bits; // @[pearray.scala 101:13]
  wire  PE_47_io_sig_stat2trans; // @[pearray.scala 101:13]
  wire  PE_48_clock; // @[pearray.scala 101:13]
  wire  PE_48_reset; // @[pearray.scala 101:13]
  wire [7:0] PE_48_io_data_2_in_bits; // @[pearray.scala 101:13]
  wire [7:0] PE_48_io_data_2_out_bits; // @[pearray.scala 101:13]
  wire  PE_48_io_data_1_in_valid; // @[pearray.scala 101:13]
  wire [7:0] PE_48_io_data_1_in_bits; // @[pearray.scala 101:13]
  wire  PE_48_io_data_1_out_valid; // @[pearray.scala 101:13]
  wire [7:0] PE_48_io_data_1_out_bits; // @[pearray.scala 101:13]
  wire  PE_48_io_data_0_in_valid; // @[pearray.scala 101:13]
  wire [7:0] PE_48_io_data_0_in_bits; // @[pearray.scala 101:13]
  wire  PE_48_io_data_0_out_valid; // @[pearray.scala 101:13]
  wire [7:0] PE_48_io_data_0_out_bits; // @[pearray.scala 101:13]
  wire  PE_48_io_sig_stat2trans; // @[pearray.scala 101:13]
  wire  PE_49_clock; // @[pearray.scala 101:13]
  wire  PE_49_reset; // @[pearray.scala 101:13]
  wire [7:0] PE_49_io_data_2_in_bits; // @[pearray.scala 101:13]
  wire [7:0] PE_49_io_data_2_out_bits; // @[pearray.scala 101:13]
  wire  PE_49_io_data_1_in_valid; // @[pearray.scala 101:13]
  wire [7:0] PE_49_io_data_1_in_bits; // @[pearray.scala 101:13]
  wire  PE_49_io_data_1_out_valid; // @[pearray.scala 101:13]
  wire [7:0] PE_49_io_data_1_out_bits; // @[pearray.scala 101:13]
  wire  PE_49_io_data_0_in_valid; // @[pearray.scala 101:13]
  wire [7:0] PE_49_io_data_0_in_bits; // @[pearray.scala 101:13]
  wire  PE_49_io_data_0_out_valid; // @[pearray.scala 101:13]
  wire [7:0] PE_49_io_data_0_out_bits; // @[pearray.scala 101:13]
  wire  PE_49_io_sig_stat2trans; // @[pearray.scala 101:13]
  wire  PE_50_clock; // @[pearray.scala 101:13]
  wire  PE_50_reset; // @[pearray.scala 101:13]
  wire [7:0] PE_50_io_data_2_in_bits; // @[pearray.scala 101:13]
  wire [7:0] PE_50_io_data_2_out_bits; // @[pearray.scala 101:13]
  wire  PE_50_io_data_1_in_valid; // @[pearray.scala 101:13]
  wire [7:0] PE_50_io_data_1_in_bits; // @[pearray.scala 101:13]
  wire  PE_50_io_data_1_out_valid; // @[pearray.scala 101:13]
  wire [7:0] PE_50_io_data_1_out_bits; // @[pearray.scala 101:13]
  wire  PE_50_io_data_0_in_valid; // @[pearray.scala 101:13]
  wire [7:0] PE_50_io_data_0_in_bits; // @[pearray.scala 101:13]
  wire  PE_50_io_data_0_out_valid; // @[pearray.scala 101:13]
  wire [7:0] PE_50_io_data_0_out_bits; // @[pearray.scala 101:13]
  wire  PE_50_io_sig_stat2trans; // @[pearray.scala 101:13]
  wire  PE_51_clock; // @[pearray.scala 101:13]
  wire  PE_51_reset; // @[pearray.scala 101:13]
  wire [7:0] PE_51_io_data_2_in_bits; // @[pearray.scala 101:13]
  wire [7:0] PE_51_io_data_2_out_bits; // @[pearray.scala 101:13]
  wire  PE_51_io_data_1_in_valid; // @[pearray.scala 101:13]
  wire [7:0] PE_51_io_data_1_in_bits; // @[pearray.scala 101:13]
  wire  PE_51_io_data_1_out_valid; // @[pearray.scala 101:13]
  wire [7:0] PE_51_io_data_1_out_bits; // @[pearray.scala 101:13]
  wire  PE_51_io_data_0_in_valid; // @[pearray.scala 101:13]
  wire [7:0] PE_51_io_data_0_in_bits; // @[pearray.scala 101:13]
  wire  PE_51_io_data_0_out_valid; // @[pearray.scala 101:13]
  wire [7:0] PE_51_io_data_0_out_bits; // @[pearray.scala 101:13]
  wire  PE_51_io_sig_stat2trans; // @[pearray.scala 101:13]
  wire  PE_52_clock; // @[pearray.scala 101:13]
  wire  PE_52_reset; // @[pearray.scala 101:13]
  wire [7:0] PE_52_io_data_2_in_bits; // @[pearray.scala 101:13]
  wire [7:0] PE_52_io_data_2_out_bits; // @[pearray.scala 101:13]
  wire  PE_52_io_data_1_in_valid; // @[pearray.scala 101:13]
  wire [7:0] PE_52_io_data_1_in_bits; // @[pearray.scala 101:13]
  wire  PE_52_io_data_1_out_valid; // @[pearray.scala 101:13]
  wire [7:0] PE_52_io_data_1_out_bits; // @[pearray.scala 101:13]
  wire  PE_52_io_data_0_in_valid; // @[pearray.scala 101:13]
  wire [7:0] PE_52_io_data_0_in_bits; // @[pearray.scala 101:13]
  wire  PE_52_io_data_0_out_valid; // @[pearray.scala 101:13]
  wire [7:0] PE_52_io_data_0_out_bits; // @[pearray.scala 101:13]
  wire  PE_52_io_sig_stat2trans; // @[pearray.scala 101:13]
  wire  PE_53_clock; // @[pearray.scala 101:13]
  wire  PE_53_reset; // @[pearray.scala 101:13]
  wire [7:0] PE_53_io_data_2_in_bits; // @[pearray.scala 101:13]
  wire [7:0] PE_53_io_data_2_out_bits; // @[pearray.scala 101:13]
  wire  PE_53_io_data_1_in_valid; // @[pearray.scala 101:13]
  wire [7:0] PE_53_io_data_1_in_bits; // @[pearray.scala 101:13]
  wire  PE_53_io_data_1_out_valid; // @[pearray.scala 101:13]
  wire [7:0] PE_53_io_data_1_out_bits; // @[pearray.scala 101:13]
  wire  PE_53_io_data_0_in_valid; // @[pearray.scala 101:13]
  wire [7:0] PE_53_io_data_0_in_bits; // @[pearray.scala 101:13]
  wire  PE_53_io_data_0_out_valid; // @[pearray.scala 101:13]
  wire [7:0] PE_53_io_data_0_out_bits; // @[pearray.scala 101:13]
  wire  PE_53_io_sig_stat2trans; // @[pearray.scala 101:13]
  wire  PE_54_clock; // @[pearray.scala 101:13]
  wire  PE_54_reset; // @[pearray.scala 101:13]
  wire [7:0] PE_54_io_data_2_in_bits; // @[pearray.scala 101:13]
  wire [7:0] PE_54_io_data_2_out_bits; // @[pearray.scala 101:13]
  wire  PE_54_io_data_1_in_valid; // @[pearray.scala 101:13]
  wire [7:0] PE_54_io_data_1_in_bits; // @[pearray.scala 101:13]
  wire  PE_54_io_data_1_out_valid; // @[pearray.scala 101:13]
  wire [7:0] PE_54_io_data_1_out_bits; // @[pearray.scala 101:13]
  wire  PE_54_io_data_0_in_valid; // @[pearray.scala 101:13]
  wire [7:0] PE_54_io_data_0_in_bits; // @[pearray.scala 101:13]
  wire  PE_54_io_data_0_out_valid; // @[pearray.scala 101:13]
  wire [7:0] PE_54_io_data_0_out_bits; // @[pearray.scala 101:13]
  wire  PE_54_io_sig_stat2trans; // @[pearray.scala 101:13]
  wire  PE_55_clock; // @[pearray.scala 101:13]
  wire  PE_55_reset; // @[pearray.scala 101:13]
  wire [7:0] PE_55_io_data_2_in_bits; // @[pearray.scala 101:13]
  wire [7:0] PE_55_io_data_2_out_bits; // @[pearray.scala 101:13]
  wire  PE_55_io_data_1_in_valid; // @[pearray.scala 101:13]
  wire [7:0] PE_55_io_data_1_in_bits; // @[pearray.scala 101:13]
  wire  PE_55_io_data_1_out_valid; // @[pearray.scala 101:13]
  wire [7:0] PE_55_io_data_1_out_bits; // @[pearray.scala 101:13]
  wire  PE_55_io_data_0_in_valid; // @[pearray.scala 101:13]
  wire [7:0] PE_55_io_data_0_in_bits; // @[pearray.scala 101:13]
  wire  PE_55_io_data_0_out_valid; // @[pearray.scala 101:13]
  wire [7:0] PE_55_io_data_0_out_bits; // @[pearray.scala 101:13]
  wire  PE_55_io_sig_stat2trans; // @[pearray.scala 101:13]
  wire  PE_56_clock; // @[pearray.scala 101:13]
  wire  PE_56_reset; // @[pearray.scala 101:13]
  wire [7:0] PE_56_io_data_2_in_bits; // @[pearray.scala 101:13]
  wire [7:0] PE_56_io_data_2_out_bits; // @[pearray.scala 101:13]
  wire  PE_56_io_data_1_in_valid; // @[pearray.scala 101:13]
  wire [7:0] PE_56_io_data_1_in_bits; // @[pearray.scala 101:13]
  wire  PE_56_io_data_1_out_valid; // @[pearray.scala 101:13]
  wire [7:0] PE_56_io_data_1_out_bits; // @[pearray.scala 101:13]
  wire  PE_56_io_data_0_in_valid; // @[pearray.scala 101:13]
  wire [7:0] PE_56_io_data_0_in_bits; // @[pearray.scala 101:13]
  wire  PE_56_io_data_0_out_valid; // @[pearray.scala 101:13]
  wire [7:0] PE_56_io_data_0_out_bits; // @[pearray.scala 101:13]
  wire  PE_56_io_sig_stat2trans; // @[pearray.scala 101:13]
  wire  PE_57_clock; // @[pearray.scala 101:13]
  wire  PE_57_reset; // @[pearray.scala 101:13]
  wire [7:0] PE_57_io_data_2_in_bits; // @[pearray.scala 101:13]
  wire [7:0] PE_57_io_data_2_out_bits; // @[pearray.scala 101:13]
  wire  PE_57_io_data_1_in_valid; // @[pearray.scala 101:13]
  wire [7:0] PE_57_io_data_1_in_bits; // @[pearray.scala 101:13]
  wire  PE_57_io_data_1_out_valid; // @[pearray.scala 101:13]
  wire [7:0] PE_57_io_data_1_out_bits; // @[pearray.scala 101:13]
  wire  PE_57_io_data_0_in_valid; // @[pearray.scala 101:13]
  wire [7:0] PE_57_io_data_0_in_bits; // @[pearray.scala 101:13]
  wire  PE_57_io_data_0_out_valid; // @[pearray.scala 101:13]
  wire [7:0] PE_57_io_data_0_out_bits; // @[pearray.scala 101:13]
  wire  PE_57_io_sig_stat2trans; // @[pearray.scala 101:13]
  wire  PE_58_clock; // @[pearray.scala 101:13]
  wire  PE_58_reset; // @[pearray.scala 101:13]
  wire [7:0] PE_58_io_data_2_in_bits; // @[pearray.scala 101:13]
  wire [7:0] PE_58_io_data_2_out_bits; // @[pearray.scala 101:13]
  wire  PE_58_io_data_1_in_valid; // @[pearray.scala 101:13]
  wire [7:0] PE_58_io_data_1_in_bits; // @[pearray.scala 101:13]
  wire  PE_58_io_data_1_out_valid; // @[pearray.scala 101:13]
  wire [7:0] PE_58_io_data_1_out_bits; // @[pearray.scala 101:13]
  wire  PE_58_io_data_0_in_valid; // @[pearray.scala 101:13]
  wire [7:0] PE_58_io_data_0_in_bits; // @[pearray.scala 101:13]
  wire  PE_58_io_data_0_out_valid; // @[pearray.scala 101:13]
  wire [7:0] PE_58_io_data_0_out_bits; // @[pearray.scala 101:13]
  wire  PE_58_io_sig_stat2trans; // @[pearray.scala 101:13]
  wire  PE_59_clock; // @[pearray.scala 101:13]
  wire  PE_59_reset; // @[pearray.scala 101:13]
  wire [7:0] PE_59_io_data_2_in_bits; // @[pearray.scala 101:13]
  wire [7:0] PE_59_io_data_2_out_bits; // @[pearray.scala 101:13]
  wire  PE_59_io_data_1_in_valid; // @[pearray.scala 101:13]
  wire [7:0] PE_59_io_data_1_in_bits; // @[pearray.scala 101:13]
  wire  PE_59_io_data_1_out_valid; // @[pearray.scala 101:13]
  wire [7:0] PE_59_io_data_1_out_bits; // @[pearray.scala 101:13]
  wire  PE_59_io_data_0_in_valid; // @[pearray.scala 101:13]
  wire [7:0] PE_59_io_data_0_in_bits; // @[pearray.scala 101:13]
  wire  PE_59_io_data_0_out_valid; // @[pearray.scala 101:13]
  wire [7:0] PE_59_io_data_0_out_bits; // @[pearray.scala 101:13]
  wire  PE_59_io_sig_stat2trans; // @[pearray.scala 101:13]
  wire  PE_60_clock; // @[pearray.scala 101:13]
  wire  PE_60_reset; // @[pearray.scala 101:13]
  wire [7:0] PE_60_io_data_2_in_bits; // @[pearray.scala 101:13]
  wire [7:0] PE_60_io_data_2_out_bits; // @[pearray.scala 101:13]
  wire  PE_60_io_data_1_in_valid; // @[pearray.scala 101:13]
  wire [7:0] PE_60_io_data_1_in_bits; // @[pearray.scala 101:13]
  wire  PE_60_io_data_1_out_valid; // @[pearray.scala 101:13]
  wire [7:0] PE_60_io_data_1_out_bits; // @[pearray.scala 101:13]
  wire  PE_60_io_data_0_in_valid; // @[pearray.scala 101:13]
  wire [7:0] PE_60_io_data_0_in_bits; // @[pearray.scala 101:13]
  wire  PE_60_io_data_0_out_valid; // @[pearray.scala 101:13]
  wire [7:0] PE_60_io_data_0_out_bits; // @[pearray.scala 101:13]
  wire  PE_60_io_sig_stat2trans; // @[pearray.scala 101:13]
  wire  PE_61_clock; // @[pearray.scala 101:13]
  wire  PE_61_reset; // @[pearray.scala 101:13]
  wire [7:0] PE_61_io_data_2_in_bits; // @[pearray.scala 101:13]
  wire [7:0] PE_61_io_data_2_out_bits; // @[pearray.scala 101:13]
  wire  PE_61_io_data_1_in_valid; // @[pearray.scala 101:13]
  wire [7:0] PE_61_io_data_1_in_bits; // @[pearray.scala 101:13]
  wire  PE_61_io_data_1_out_valid; // @[pearray.scala 101:13]
  wire [7:0] PE_61_io_data_1_out_bits; // @[pearray.scala 101:13]
  wire  PE_61_io_data_0_in_valid; // @[pearray.scala 101:13]
  wire [7:0] PE_61_io_data_0_in_bits; // @[pearray.scala 101:13]
  wire  PE_61_io_data_0_out_valid; // @[pearray.scala 101:13]
  wire [7:0] PE_61_io_data_0_out_bits; // @[pearray.scala 101:13]
  wire  PE_61_io_sig_stat2trans; // @[pearray.scala 101:13]
  wire  PE_62_clock; // @[pearray.scala 101:13]
  wire  PE_62_reset; // @[pearray.scala 101:13]
  wire [7:0] PE_62_io_data_2_in_bits; // @[pearray.scala 101:13]
  wire [7:0] PE_62_io_data_2_out_bits; // @[pearray.scala 101:13]
  wire  PE_62_io_data_1_in_valid; // @[pearray.scala 101:13]
  wire [7:0] PE_62_io_data_1_in_bits; // @[pearray.scala 101:13]
  wire  PE_62_io_data_1_out_valid; // @[pearray.scala 101:13]
  wire [7:0] PE_62_io_data_1_out_bits; // @[pearray.scala 101:13]
  wire  PE_62_io_data_0_in_valid; // @[pearray.scala 101:13]
  wire [7:0] PE_62_io_data_0_in_bits; // @[pearray.scala 101:13]
  wire  PE_62_io_data_0_out_valid; // @[pearray.scala 101:13]
  wire [7:0] PE_62_io_data_0_out_bits; // @[pearray.scala 101:13]
  wire  PE_62_io_sig_stat2trans; // @[pearray.scala 101:13]
  wire  PE_63_clock; // @[pearray.scala 101:13]
  wire  PE_63_reset; // @[pearray.scala 101:13]
  wire [7:0] PE_63_io_data_2_in_bits; // @[pearray.scala 101:13]
  wire [7:0] PE_63_io_data_2_out_bits; // @[pearray.scala 101:13]
  wire  PE_63_io_data_1_in_valid; // @[pearray.scala 101:13]
  wire [7:0] PE_63_io_data_1_in_bits; // @[pearray.scala 101:13]
  wire  PE_63_io_data_1_out_valid; // @[pearray.scala 101:13]
  wire [7:0] PE_63_io_data_1_out_bits; // @[pearray.scala 101:13]
  wire  PE_63_io_data_0_in_valid; // @[pearray.scala 101:13]
  wire [7:0] PE_63_io_data_0_in_bits; // @[pearray.scala 101:13]
  wire  PE_63_io_data_0_out_valid; // @[pearray.scala 101:13]
  wire [7:0] PE_63_io_data_0_out_bits; // @[pearray.scala 101:13]
  wire  PE_63_io_sig_stat2trans; // @[pearray.scala 101:13]
  wire  PE_64_clock; // @[pearray.scala 101:13]
  wire  PE_64_reset; // @[pearray.scala 101:13]
  wire [7:0] PE_64_io_data_2_in_bits; // @[pearray.scala 101:13]
  wire [7:0] PE_64_io_data_2_out_bits; // @[pearray.scala 101:13]
  wire  PE_64_io_data_1_in_valid; // @[pearray.scala 101:13]
  wire [7:0] PE_64_io_data_1_in_bits; // @[pearray.scala 101:13]
  wire  PE_64_io_data_1_out_valid; // @[pearray.scala 101:13]
  wire [7:0] PE_64_io_data_1_out_bits; // @[pearray.scala 101:13]
  wire  PE_64_io_data_0_in_valid; // @[pearray.scala 101:13]
  wire [7:0] PE_64_io_data_0_in_bits; // @[pearray.scala 101:13]
  wire  PE_64_io_data_0_out_valid; // @[pearray.scala 101:13]
  wire [7:0] PE_64_io_data_0_out_bits; // @[pearray.scala 101:13]
  wire  PE_64_io_sig_stat2trans; // @[pearray.scala 101:13]
  wire  PE_65_clock; // @[pearray.scala 101:13]
  wire  PE_65_reset; // @[pearray.scala 101:13]
  wire [7:0] PE_65_io_data_2_in_bits; // @[pearray.scala 101:13]
  wire [7:0] PE_65_io_data_2_out_bits; // @[pearray.scala 101:13]
  wire  PE_65_io_data_1_in_valid; // @[pearray.scala 101:13]
  wire [7:0] PE_65_io_data_1_in_bits; // @[pearray.scala 101:13]
  wire  PE_65_io_data_1_out_valid; // @[pearray.scala 101:13]
  wire [7:0] PE_65_io_data_1_out_bits; // @[pearray.scala 101:13]
  wire  PE_65_io_data_0_in_valid; // @[pearray.scala 101:13]
  wire [7:0] PE_65_io_data_0_in_bits; // @[pearray.scala 101:13]
  wire  PE_65_io_data_0_out_valid; // @[pearray.scala 101:13]
  wire [7:0] PE_65_io_data_0_out_bits; // @[pearray.scala 101:13]
  wire  PE_65_io_sig_stat2trans; // @[pearray.scala 101:13]
  wire  PE_66_clock; // @[pearray.scala 101:13]
  wire  PE_66_reset; // @[pearray.scala 101:13]
  wire [7:0] PE_66_io_data_2_in_bits; // @[pearray.scala 101:13]
  wire [7:0] PE_66_io_data_2_out_bits; // @[pearray.scala 101:13]
  wire  PE_66_io_data_1_in_valid; // @[pearray.scala 101:13]
  wire [7:0] PE_66_io_data_1_in_bits; // @[pearray.scala 101:13]
  wire  PE_66_io_data_1_out_valid; // @[pearray.scala 101:13]
  wire [7:0] PE_66_io_data_1_out_bits; // @[pearray.scala 101:13]
  wire  PE_66_io_data_0_in_valid; // @[pearray.scala 101:13]
  wire [7:0] PE_66_io_data_0_in_bits; // @[pearray.scala 101:13]
  wire  PE_66_io_data_0_out_valid; // @[pearray.scala 101:13]
  wire [7:0] PE_66_io_data_0_out_bits; // @[pearray.scala 101:13]
  wire  PE_66_io_sig_stat2trans; // @[pearray.scala 101:13]
  wire  PE_67_clock; // @[pearray.scala 101:13]
  wire  PE_67_reset; // @[pearray.scala 101:13]
  wire [7:0] PE_67_io_data_2_in_bits; // @[pearray.scala 101:13]
  wire [7:0] PE_67_io_data_2_out_bits; // @[pearray.scala 101:13]
  wire  PE_67_io_data_1_in_valid; // @[pearray.scala 101:13]
  wire [7:0] PE_67_io_data_1_in_bits; // @[pearray.scala 101:13]
  wire  PE_67_io_data_1_out_valid; // @[pearray.scala 101:13]
  wire [7:0] PE_67_io_data_1_out_bits; // @[pearray.scala 101:13]
  wire  PE_67_io_data_0_in_valid; // @[pearray.scala 101:13]
  wire [7:0] PE_67_io_data_0_in_bits; // @[pearray.scala 101:13]
  wire  PE_67_io_data_0_out_valid; // @[pearray.scala 101:13]
  wire [7:0] PE_67_io_data_0_out_bits; // @[pearray.scala 101:13]
  wire  PE_67_io_sig_stat2trans; // @[pearray.scala 101:13]
  wire  PE_68_clock; // @[pearray.scala 101:13]
  wire  PE_68_reset; // @[pearray.scala 101:13]
  wire [7:0] PE_68_io_data_2_in_bits; // @[pearray.scala 101:13]
  wire [7:0] PE_68_io_data_2_out_bits; // @[pearray.scala 101:13]
  wire  PE_68_io_data_1_in_valid; // @[pearray.scala 101:13]
  wire [7:0] PE_68_io_data_1_in_bits; // @[pearray.scala 101:13]
  wire  PE_68_io_data_1_out_valid; // @[pearray.scala 101:13]
  wire [7:0] PE_68_io_data_1_out_bits; // @[pearray.scala 101:13]
  wire  PE_68_io_data_0_in_valid; // @[pearray.scala 101:13]
  wire [7:0] PE_68_io_data_0_in_bits; // @[pearray.scala 101:13]
  wire  PE_68_io_data_0_out_valid; // @[pearray.scala 101:13]
  wire [7:0] PE_68_io_data_0_out_bits; // @[pearray.scala 101:13]
  wire  PE_68_io_sig_stat2trans; // @[pearray.scala 101:13]
  wire  PE_69_clock; // @[pearray.scala 101:13]
  wire  PE_69_reset; // @[pearray.scala 101:13]
  wire [7:0] PE_69_io_data_2_in_bits; // @[pearray.scala 101:13]
  wire [7:0] PE_69_io_data_2_out_bits; // @[pearray.scala 101:13]
  wire  PE_69_io_data_1_in_valid; // @[pearray.scala 101:13]
  wire [7:0] PE_69_io_data_1_in_bits; // @[pearray.scala 101:13]
  wire  PE_69_io_data_1_out_valid; // @[pearray.scala 101:13]
  wire [7:0] PE_69_io_data_1_out_bits; // @[pearray.scala 101:13]
  wire  PE_69_io_data_0_in_valid; // @[pearray.scala 101:13]
  wire [7:0] PE_69_io_data_0_in_bits; // @[pearray.scala 101:13]
  wire  PE_69_io_data_0_out_valid; // @[pearray.scala 101:13]
  wire [7:0] PE_69_io_data_0_out_bits; // @[pearray.scala 101:13]
  wire  PE_69_io_sig_stat2trans; // @[pearray.scala 101:13]
  wire  PE_70_clock; // @[pearray.scala 101:13]
  wire  PE_70_reset; // @[pearray.scala 101:13]
  wire [7:0] PE_70_io_data_2_in_bits; // @[pearray.scala 101:13]
  wire [7:0] PE_70_io_data_2_out_bits; // @[pearray.scala 101:13]
  wire  PE_70_io_data_1_in_valid; // @[pearray.scala 101:13]
  wire [7:0] PE_70_io_data_1_in_bits; // @[pearray.scala 101:13]
  wire  PE_70_io_data_1_out_valid; // @[pearray.scala 101:13]
  wire [7:0] PE_70_io_data_1_out_bits; // @[pearray.scala 101:13]
  wire  PE_70_io_data_0_in_valid; // @[pearray.scala 101:13]
  wire [7:0] PE_70_io_data_0_in_bits; // @[pearray.scala 101:13]
  wire  PE_70_io_data_0_out_valid; // @[pearray.scala 101:13]
  wire [7:0] PE_70_io_data_0_out_bits; // @[pearray.scala 101:13]
  wire  PE_70_io_sig_stat2trans; // @[pearray.scala 101:13]
  wire  PE_71_clock; // @[pearray.scala 101:13]
  wire  PE_71_reset; // @[pearray.scala 101:13]
  wire [7:0] PE_71_io_data_2_in_bits; // @[pearray.scala 101:13]
  wire [7:0] PE_71_io_data_2_out_bits; // @[pearray.scala 101:13]
  wire  PE_71_io_data_1_in_valid; // @[pearray.scala 101:13]
  wire [7:0] PE_71_io_data_1_in_bits; // @[pearray.scala 101:13]
  wire  PE_71_io_data_1_out_valid; // @[pearray.scala 101:13]
  wire [7:0] PE_71_io_data_1_out_bits; // @[pearray.scala 101:13]
  wire  PE_71_io_data_0_in_valid; // @[pearray.scala 101:13]
  wire [7:0] PE_71_io_data_0_in_bits; // @[pearray.scala 101:13]
  wire  PE_71_io_data_0_out_valid; // @[pearray.scala 101:13]
  wire [7:0] PE_71_io_data_0_out_bits; // @[pearray.scala 101:13]
  wire  PE_71_io_sig_stat2trans; // @[pearray.scala 101:13]
  wire  PE_72_clock; // @[pearray.scala 101:13]
  wire  PE_72_reset; // @[pearray.scala 101:13]
  wire [7:0] PE_72_io_data_2_in_bits; // @[pearray.scala 101:13]
  wire [7:0] PE_72_io_data_2_out_bits; // @[pearray.scala 101:13]
  wire  PE_72_io_data_1_in_valid; // @[pearray.scala 101:13]
  wire [7:0] PE_72_io_data_1_in_bits; // @[pearray.scala 101:13]
  wire  PE_72_io_data_1_out_valid; // @[pearray.scala 101:13]
  wire [7:0] PE_72_io_data_1_out_bits; // @[pearray.scala 101:13]
  wire  PE_72_io_data_0_in_valid; // @[pearray.scala 101:13]
  wire [7:0] PE_72_io_data_0_in_bits; // @[pearray.scala 101:13]
  wire  PE_72_io_data_0_out_valid; // @[pearray.scala 101:13]
  wire [7:0] PE_72_io_data_0_out_bits; // @[pearray.scala 101:13]
  wire  PE_72_io_sig_stat2trans; // @[pearray.scala 101:13]
  wire  PE_73_clock; // @[pearray.scala 101:13]
  wire  PE_73_reset; // @[pearray.scala 101:13]
  wire [7:0] PE_73_io_data_2_in_bits; // @[pearray.scala 101:13]
  wire [7:0] PE_73_io_data_2_out_bits; // @[pearray.scala 101:13]
  wire  PE_73_io_data_1_in_valid; // @[pearray.scala 101:13]
  wire [7:0] PE_73_io_data_1_in_bits; // @[pearray.scala 101:13]
  wire  PE_73_io_data_1_out_valid; // @[pearray.scala 101:13]
  wire [7:0] PE_73_io_data_1_out_bits; // @[pearray.scala 101:13]
  wire  PE_73_io_data_0_in_valid; // @[pearray.scala 101:13]
  wire [7:0] PE_73_io_data_0_in_bits; // @[pearray.scala 101:13]
  wire  PE_73_io_data_0_out_valid; // @[pearray.scala 101:13]
  wire [7:0] PE_73_io_data_0_out_bits; // @[pearray.scala 101:13]
  wire  PE_73_io_sig_stat2trans; // @[pearray.scala 101:13]
  wire  PE_74_clock; // @[pearray.scala 101:13]
  wire  PE_74_reset; // @[pearray.scala 101:13]
  wire [7:0] PE_74_io_data_2_in_bits; // @[pearray.scala 101:13]
  wire [7:0] PE_74_io_data_2_out_bits; // @[pearray.scala 101:13]
  wire  PE_74_io_data_1_in_valid; // @[pearray.scala 101:13]
  wire [7:0] PE_74_io_data_1_in_bits; // @[pearray.scala 101:13]
  wire  PE_74_io_data_1_out_valid; // @[pearray.scala 101:13]
  wire [7:0] PE_74_io_data_1_out_bits; // @[pearray.scala 101:13]
  wire  PE_74_io_data_0_in_valid; // @[pearray.scala 101:13]
  wire [7:0] PE_74_io_data_0_in_bits; // @[pearray.scala 101:13]
  wire  PE_74_io_data_0_out_valid; // @[pearray.scala 101:13]
  wire [7:0] PE_74_io_data_0_out_bits; // @[pearray.scala 101:13]
  wire  PE_74_io_sig_stat2trans; // @[pearray.scala 101:13]
  wire  PE_75_clock; // @[pearray.scala 101:13]
  wire  PE_75_reset; // @[pearray.scala 101:13]
  wire [7:0] PE_75_io_data_2_in_bits; // @[pearray.scala 101:13]
  wire [7:0] PE_75_io_data_2_out_bits; // @[pearray.scala 101:13]
  wire  PE_75_io_data_1_in_valid; // @[pearray.scala 101:13]
  wire [7:0] PE_75_io_data_1_in_bits; // @[pearray.scala 101:13]
  wire  PE_75_io_data_1_out_valid; // @[pearray.scala 101:13]
  wire [7:0] PE_75_io_data_1_out_bits; // @[pearray.scala 101:13]
  wire  PE_75_io_data_0_in_valid; // @[pearray.scala 101:13]
  wire [7:0] PE_75_io_data_0_in_bits; // @[pearray.scala 101:13]
  wire  PE_75_io_data_0_out_valid; // @[pearray.scala 101:13]
  wire [7:0] PE_75_io_data_0_out_bits; // @[pearray.scala 101:13]
  wire  PE_75_io_sig_stat2trans; // @[pearray.scala 101:13]
  wire  PE_76_clock; // @[pearray.scala 101:13]
  wire  PE_76_reset; // @[pearray.scala 101:13]
  wire [7:0] PE_76_io_data_2_in_bits; // @[pearray.scala 101:13]
  wire [7:0] PE_76_io_data_2_out_bits; // @[pearray.scala 101:13]
  wire  PE_76_io_data_1_in_valid; // @[pearray.scala 101:13]
  wire [7:0] PE_76_io_data_1_in_bits; // @[pearray.scala 101:13]
  wire  PE_76_io_data_1_out_valid; // @[pearray.scala 101:13]
  wire [7:0] PE_76_io_data_1_out_bits; // @[pearray.scala 101:13]
  wire  PE_76_io_data_0_in_valid; // @[pearray.scala 101:13]
  wire [7:0] PE_76_io_data_0_in_bits; // @[pearray.scala 101:13]
  wire  PE_76_io_data_0_out_valid; // @[pearray.scala 101:13]
  wire [7:0] PE_76_io_data_0_out_bits; // @[pearray.scala 101:13]
  wire  PE_76_io_sig_stat2trans; // @[pearray.scala 101:13]
  wire  PE_77_clock; // @[pearray.scala 101:13]
  wire  PE_77_reset; // @[pearray.scala 101:13]
  wire [7:0] PE_77_io_data_2_in_bits; // @[pearray.scala 101:13]
  wire [7:0] PE_77_io_data_2_out_bits; // @[pearray.scala 101:13]
  wire  PE_77_io_data_1_in_valid; // @[pearray.scala 101:13]
  wire [7:0] PE_77_io_data_1_in_bits; // @[pearray.scala 101:13]
  wire  PE_77_io_data_1_out_valid; // @[pearray.scala 101:13]
  wire [7:0] PE_77_io_data_1_out_bits; // @[pearray.scala 101:13]
  wire  PE_77_io_data_0_in_valid; // @[pearray.scala 101:13]
  wire [7:0] PE_77_io_data_0_in_bits; // @[pearray.scala 101:13]
  wire  PE_77_io_data_0_out_valid; // @[pearray.scala 101:13]
  wire [7:0] PE_77_io_data_0_out_bits; // @[pearray.scala 101:13]
  wire  PE_77_io_sig_stat2trans; // @[pearray.scala 101:13]
  wire  PE_78_clock; // @[pearray.scala 101:13]
  wire  PE_78_reset; // @[pearray.scala 101:13]
  wire [7:0] PE_78_io_data_2_in_bits; // @[pearray.scala 101:13]
  wire [7:0] PE_78_io_data_2_out_bits; // @[pearray.scala 101:13]
  wire  PE_78_io_data_1_in_valid; // @[pearray.scala 101:13]
  wire [7:0] PE_78_io_data_1_in_bits; // @[pearray.scala 101:13]
  wire  PE_78_io_data_1_out_valid; // @[pearray.scala 101:13]
  wire [7:0] PE_78_io_data_1_out_bits; // @[pearray.scala 101:13]
  wire  PE_78_io_data_0_in_valid; // @[pearray.scala 101:13]
  wire [7:0] PE_78_io_data_0_in_bits; // @[pearray.scala 101:13]
  wire  PE_78_io_data_0_out_valid; // @[pearray.scala 101:13]
  wire [7:0] PE_78_io_data_0_out_bits; // @[pearray.scala 101:13]
  wire  PE_78_io_sig_stat2trans; // @[pearray.scala 101:13]
  wire  PE_79_clock; // @[pearray.scala 101:13]
  wire  PE_79_reset; // @[pearray.scala 101:13]
  wire [7:0] PE_79_io_data_2_in_bits; // @[pearray.scala 101:13]
  wire [7:0] PE_79_io_data_2_out_bits; // @[pearray.scala 101:13]
  wire  PE_79_io_data_1_in_valid; // @[pearray.scala 101:13]
  wire [7:0] PE_79_io_data_1_in_bits; // @[pearray.scala 101:13]
  wire  PE_79_io_data_1_out_valid; // @[pearray.scala 101:13]
  wire [7:0] PE_79_io_data_1_out_bits; // @[pearray.scala 101:13]
  wire  PE_79_io_data_0_in_valid; // @[pearray.scala 101:13]
  wire [7:0] PE_79_io_data_0_in_bits; // @[pearray.scala 101:13]
  wire  PE_79_io_data_0_out_valid; // @[pearray.scala 101:13]
  wire [7:0] PE_79_io_data_0_out_bits; // @[pearray.scala 101:13]
  wire  PE_79_io_sig_stat2trans; // @[pearray.scala 101:13]
  wire  PE_80_clock; // @[pearray.scala 101:13]
  wire  PE_80_reset; // @[pearray.scala 101:13]
  wire [7:0] PE_80_io_data_2_in_bits; // @[pearray.scala 101:13]
  wire [7:0] PE_80_io_data_2_out_bits; // @[pearray.scala 101:13]
  wire  PE_80_io_data_1_in_valid; // @[pearray.scala 101:13]
  wire [7:0] PE_80_io_data_1_in_bits; // @[pearray.scala 101:13]
  wire  PE_80_io_data_1_out_valid; // @[pearray.scala 101:13]
  wire [7:0] PE_80_io_data_1_out_bits; // @[pearray.scala 101:13]
  wire  PE_80_io_data_0_in_valid; // @[pearray.scala 101:13]
  wire [7:0] PE_80_io_data_0_in_bits; // @[pearray.scala 101:13]
  wire  PE_80_io_data_0_out_valid; // @[pearray.scala 101:13]
  wire [7:0] PE_80_io_data_0_out_bits; // @[pearray.scala 101:13]
  wire  PE_80_io_sig_stat2trans; // @[pearray.scala 101:13]
  wire  PE_81_clock; // @[pearray.scala 101:13]
  wire  PE_81_reset; // @[pearray.scala 101:13]
  wire [7:0] PE_81_io_data_2_in_bits; // @[pearray.scala 101:13]
  wire [7:0] PE_81_io_data_2_out_bits; // @[pearray.scala 101:13]
  wire  PE_81_io_data_1_in_valid; // @[pearray.scala 101:13]
  wire [7:0] PE_81_io_data_1_in_bits; // @[pearray.scala 101:13]
  wire  PE_81_io_data_1_out_valid; // @[pearray.scala 101:13]
  wire [7:0] PE_81_io_data_1_out_bits; // @[pearray.scala 101:13]
  wire  PE_81_io_data_0_in_valid; // @[pearray.scala 101:13]
  wire [7:0] PE_81_io_data_0_in_bits; // @[pearray.scala 101:13]
  wire  PE_81_io_data_0_out_valid; // @[pearray.scala 101:13]
  wire [7:0] PE_81_io_data_0_out_bits; // @[pearray.scala 101:13]
  wire  PE_81_io_sig_stat2trans; // @[pearray.scala 101:13]
  wire  PE_82_clock; // @[pearray.scala 101:13]
  wire  PE_82_reset; // @[pearray.scala 101:13]
  wire [7:0] PE_82_io_data_2_in_bits; // @[pearray.scala 101:13]
  wire [7:0] PE_82_io_data_2_out_bits; // @[pearray.scala 101:13]
  wire  PE_82_io_data_1_in_valid; // @[pearray.scala 101:13]
  wire [7:0] PE_82_io_data_1_in_bits; // @[pearray.scala 101:13]
  wire  PE_82_io_data_1_out_valid; // @[pearray.scala 101:13]
  wire [7:0] PE_82_io_data_1_out_bits; // @[pearray.scala 101:13]
  wire  PE_82_io_data_0_in_valid; // @[pearray.scala 101:13]
  wire [7:0] PE_82_io_data_0_in_bits; // @[pearray.scala 101:13]
  wire  PE_82_io_data_0_out_valid; // @[pearray.scala 101:13]
  wire [7:0] PE_82_io_data_0_out_bits; // @[pearray.scala 101:13]
  wire  PE_82_io_sig_stat2trans; // @[pearray.scala 101:13]
  wire  PE_83_clock; // @[pearray.scala 101:13]
  wire  PE_83_reset; // @[pearray.scala 101:13]
  wire [7:0] PE_83_io_data_2_in_bits; // @[pearray.scala 101:13]
  wire [7:0] PE_83_io_data_2_out_bits; // @[pearray.scala 101:13]
  wire  PE_83_io_data_1_in_valid; // @[pearray.scala 101:13]
  wire [7:0] PE_83_io_data_1_in_bits; // @[pearray.scala 101:13]
  wire  PE_83_io_data_1_out_valid; // @[pearray.scala 101:13]
  wire [7:0] PE_83_io_data_1_out_bits; // @[pearray.scala 101:13]
  wire  PE_83_io_data_0_in_valid; // @[pearray.scala 101:13]
  wire [7:0] PE_83_io_data_0_in_bits; // @[pearray.scala 101:13]
  wire  PE_83_io_data_0_out_valid; // @[pearray.scala 101:13]
  wire [7:0] PE_83_io_data_0_out_bits; // @[pearray.scala 101:13]
  wire  PE_83_io_sig_stat2trans; // @[pearray.scala 101:13]
  wire  PE_84_clock; // @[pearray.scala 101:13]
  wire  PE_84_reset; // @[pearray.scala 101:13]
  wire [7:0] PE_84_io_data_2_in_bits; // @[pearray.scala 101:13]
  wire [7:0] PE_84_io_data_2_out_bits; // @[pearray.scala 101:13]
  wire  PE_84_io_data_1_in_valid; // @[pearray.scala 101:13]
  wire [7:0] PE_84_io_data_1_in_bits; // @[pearray.scala 101:13]
  wire  PE_84_io_data_1_out_valid; // @[pearray.scala 101:13]
  wire [7:0] PE_84_io_data_1_out_bits; // @[pearray.scala 101:13]
  wire  PE_84_io_data_0_in_valid; // @[pearray.scala 101:13]
  wire [7:0] PE_84_io_data_0_in_bits; // @[pearray.scala 101:13]
  wire  PE_84_io_data_0_out_valid; // @[pearray.scala 101:13]
  wire [7:0] PE_84_io_data_0_out_bits; // @[pearray.scala 101:13]
  wire  PE_84_io_sig_stat2trans; // @[pearray.scala 101:13]
  wire  PE_85_clock; // @[pearray.scala 101:13]
  wire  PE_85_reset; // @[pearray.scala 101:13]
  wire [7:0] PE_85_io_data_2_in_bits; // @[pearray.scala 101:13]
  wire [7:0] PE_85_io_data_2_out_bits; // @[pearray.scala 101:13]
  wire  PE_85_io_data_1_in_valid; // @[pearray.scala 101:13]
  wire [7:0] PE_85_io_data_1_in_bits; // @[pearray.scala 101:13]
  wire  PE_85_io_data_1_out_valid; // @[pearray.scala 101:13]
  wire [7:0] PE_85_io_data_1_out_bits; // @[pearray.scala 101:13]
  wire  PE_85_io_data_0_in_valid; // @[pearray.scala 101:13]
  wire [7:0] PE_85_io_data_0_in_bits; // @[pearray.scala 101:13]
  wire  PE_85_io_data_0_out_valid; // @[pearray.scala 101:13]
  wire [7:0] PE_85_io_data_0_out_bits; // @[pearray.scala 101:13]
  wire  PE_85_io_sig_stat2trans; // @[pearray.scala 101:13]
  wire  PE_86_clock; // @[pearray.scala 101:13]
  wire  PE_86_reset; // @[pearray.scala 101:13]
  wire [7:0] PE_86_io_data_2_in_bits; // @[pearray.scala 101:13]
  wire [7:0] PE_86_io_data_2_out_bits; // @[pearray.scala 101:13]
  wire  PE_86_io_data_1_in_valid; // @[pearray.scala 101:13]
  wire [7:0] PE_86_io_data_1_in_bits; // @[pearray.scala 101:13]
  wire  PE_86_io_data_1_out_valid; // @[pearray.scala 101:13]
  wire [7:0] PE_86_io_data_1_out_bits; // @[pearray.scala 101:13]
  wire  PE_86_io_data_0_in_valid; // @[pearray.scala 101:13]
  wire [7:0] PE_86_io_data_0_in_bits; // @[pearray.scala 101:13]
  wire  PE_86_io_data_0_out_valid; // @[pearray.scala 101:13]
  wire [7:0] PE_86_io_data_0_out_bits; // @[pearray.scala 101:13]
  wire  PE_86_io_sig_stat2trans; // @[pearray.scala 101:13]
  wire  PE_87_clock; // @[pearray.scala 101:13]
  wire  PE_87_reset; // @[pearray.scala 101:13]
  wire [7:0] PE_87_io_data_2_in_bits; // @[pearray.scala 101:13]
  wire [7:0] PE_87_io_data_2_out_bits; // @[pearray.scala 101:13]
  wire  PE_87_io_data_1_in_valid; // @[pearray.scala 101:13]
  wire [7:0] PE_87_io_data_1_in_bits; // @[pearray.scala 101:13]
  wire  PE_87_io_data_1_out_valid; // @[pearray.scala 101:13]
  wire [7:0] PE_87_io_data_1_out_bits; // @[pearray.scala 101:13]
  wire  PE_87_io_data_0_in_valid; // @[pearray.scala 101:13]
  wire [7:0] PE_87_io_data_0_in_bits; // @[pearray.scala 101:13]
  wire  PE_87_io_data_0_out_valid; // @[pearray.scala 101:13]
  wire [7:0] PE_87_io_data_0_out_bits; // @[pearray.scala 101:13]
  wire  PE_87_io_sig_stat2trans; // @[pearray.scala 101:13]
  wire  PE_88_clock; // @[pearray.scala 101:13]
  wire  PE_88_reset; // @[pearray.scala 101:13]
  wire [7:0] PE_88_io_data_2_in_bits; // @[pearray.scala 101:13]
  wire [7:0] PE_88_io_data_2_out_bits; // @[pearray.scala 101:13]
  wire  PE_88_io_data_1_in_valid; // @[pearray.scala 101:13]
  wire [7:0] PE_88_io_data_1_in_bits; // @[pearray.scala 101:13]
  wire  PE_88_io_data_1_out_valid; // @[pearray.scala 101:13]
  wire [7:0] PE_88_io_data_1_out_bits; // @[pearray.scala 101:13]
  wire  PE_88_io_data_0_in_valid; // @[pearray.scala 101:13]
  wire [7:0] PE_88_io_data_0_in_bits; // @[pearray.scala 101:13]
  wire  PE_88_io_data_0_out_valid; // @[pearray.scala 101:13]
  wire [7:0] PE_88_io_data_0_out_bits; // @[pearray.scala 101:13]
  wire  PE_88_io_sig_stat2trans; // @[pearray.scala 101:13]
  wire  PE_89_clock; // @[pearray.scala 101:13]
  wire  PE_89_reset; // @[pearray.scala 101:13]
  wire [7:0] PE_89_io_data_2_in_bits; // @[pearray.scala 101:13]
  wire [7:0] PE_89_io_data_2_out_bits; // @[pearray.scala 101:13]
  wire  PE_89_io_data_1_in_valid; // @[pearray.scala 101:13]
  wire [7:0] PE_89_io_data_1_in_bits; // @[pearray.scala 101:13]
  wire  PE_89_io_data_1_out_valid; // @[pearray.scala 101:13]
  wire [7:0] PE_89_io_data_1_out_bits; // @[pearray.scala 101:13]
  wire  PE_89_io_data_0_in_valid; // @[pearray.scala 101:13]
  wire [7:0] PE_89_io_data_0_in_bits; // @[pearray.scala 101:13]
  wire  PE_89_io_data_0_out_valid; // @[pearray.scala 101:13]
  wire [7:0] PE_89_io_data_0_out_bits; // @[pearray.scala 101:13]
  wire  PE_89_io_sig_stat2trans; // @[pearray.scala 101:13]
  wire  PE_90_clock; // @[pearray.scala 101:13]
  wire  PE_90_reset; // @[pearray.scala 101:13]
  wire [7:0] PE_90_io_data_2_in_bits; // @[pearray.scala 101:13]
  wire [7:0] PE_90_io_data_2_out_bits; // @[pearray.scala 101:13]
  wire  PE_90_io_data_1_in_valid; // @[pearray.scala 101:13]
  wire [7:0] PE_90_io_data_1_in_bits; // @[pearray.scala 101:13]
  wire  PE_90_io_data_1_out_valid; // @[pearray.scala 101:13]
  wire [7:0] PE_90_io_data_1_out_bits; // @[pearray.scala 101:13]
  wire  PE_90_io_data_0_in_valid; // @[pearray.scala 101:13]
  wire [7:0] PE_90_io_data_0_in_bits; // @[pearray.scala 101:13]
  wire  PE_90_io_data_0_out_valid; // @[pearray.scala 101:13]
  wire [7:0] PE_90_io_data_0_out_bits; // @[pearray.scala 101:13]
  wire  PE_90_io_sig_stat2trans; // @[pearray.scala 101:13]
  wire  PE_91_clock; // @[pearray.scala 101:13]
  wire  PE_91_reset; // @[pearray.scala 101:13]
  wire [7:0] PE_91_io_data_2_in_bits; // @[pearray.scala 101:13]
  wire [7:0] PE_91_io_data_2_out_bits; // @[pearray.scala 101:13]
  wire  PE_91_io_data_1_in_valid; // @[pearray.scala 101:13]
  wire [7:0] PE_91_io_data_1_in_bits; // @[pearray.scala 101:13]
  wire  PE_91_io_data_1_out_valid; // @[pearray.scala 101:13]
  wire [7:0] PE_91_io_data_1_out_bits; // @[pearray.scala 101:13]
  wire  PE_91_io_data_0_in_valid; // @[pearray.scala 101:13]
  wire [7:0] PE_91_io_data_0_in_bits; // @[pearray.scala 101:13]
  wire  PE_91_io_data_0_out_valid; // @[pearray.scala 101:13]
  wire [7:0] PE_91_io_data_0_out_bits; // @[pearray.scala 101:13]
  wire  PE_91_io_sig_stat2trans; // @[pearray.scala 101:13]
  wire  PE_92_clock; // @[pearray.scala 101:13]
  wire  PE_92_reset; // @[pearray.scala 101:13]
  wire [7:0] PE_92_io_data_2_in_bits; // @[pearray.scala 101:13]
  wire [7:0] PE_92_io_data_2_out_bits; // @[pearray.scala 101:13]
  wire  PE_92_io_data_1_in_valid; // @[pearray.scala 101:13]
  wire [7:0] PE_92_io_data_1_in_bits; // @[pearray.scala 101:13]
  wire  PE_92_io_data_1_out_valid; // @[pearray.scala 101:13]
  wire [7:0] PE_92_io_data_1_out_bits; // @[pearray.scala 101:13]
  wire  PE_92_io_data_0_in_valid; // @[pearray.scala 101:13]
  wire [7:0] PE_92_io_data_0_in_bits; // @[pearray.scala 101:13]
  wire  PE_92_io_data_0_out_valid; // @[pearray.scala 101:13]
  wire [7:0] PE_92_io_data_0_out_bits; // @[pearray.scala 101:13]
  wire  PE_92_io_sig_stat2trans; // @[pearray.scala 101:13]
  wire  PE_93_clock; // @[pearray.scala 101:13]
  wire  PE_93_reset; // @[pearray.scala 101:13]
  wire [7:0] PE_93_io_data_2_in_bits; // @[pearray.scala 101:13]
  wire [7:0] PE_93_io_data_2_out_bits; // @[pearray.scala 101:13]
  wire  PE_93_io_data_1_in_valid; // @[pearray.scala 101:13]
  wire [7:0] PE_93_io_data_1_in_bits; // @[pearray.scala 101:13]
  wire  PE_93_io_data_1_out_valid; // @[pearray.scala 101:13]
  wire [7:0] PE_93_io_data_1_out_bits; // @[pearray.scala 101:13]
  wire  PE_93_io_data_0_in_valid; // @[pearray.scala 101:13]
  wire [7:0] PE_93_io_data_0_in_bits; // @[pearray.scala 101:13]
  wire  PE_93_io_data_0_out_valid; // @[pearray.scala 101:13]
  wire [7:0] PE_93_io_data_0_out_bits; // @[pearray.scala 101:13]
  wire  PE_93_io_sig_stat2trans; // @[pearray.scala 101:13]
  wire  PE_94_clock; // @[pearray.scala 101:13]
  wire  PE_94_reset; // @[pearray.scala 101:13]
  wire [7:0] PE_94_io_data_2_in_bits; // @[pearray.scala 101:13]
  wire [7:0] PE_94_io_data_2_out_bits; // @[pearray.scala 101:13]
  wire  PE_94_io_data_1_in_valid; // @[pearray.scala 101:13]
  wire [7:0] PE_94_io_data_1_in_bits; // @[pearray.scala 101:13]
  wire  PE_94_io_data_1_out_valid; // @[pearray.scala 101:13]
  wire [7:0] PE_94_io_data_1_out_bits; // @[pearray.scala 101:13]
  wire  PE_94_io_data_0_in_valid; // @[pearray.scala 101:13]
  wire [7:0] PE_94_io_data_0_in_bits; // @[pearray.scala 101:13]
  wire  PE_94_io_data_0_out_valid; // @[pearray.scala 101:13]
  wire [7:0] PE_94_io_data_0_out_bits; // @[pearray.scala 101:13]
  wire  PE_94_io_sig_stat2trans; // @[pearray.scala 101:13]
  wire  PE_95_clock; // @[pearray.scala 101:13]
  wire  PE_95_reset; // @[pearray.scala 101:13]
  wire [7:0] PE_95_io_data_2_in_bits; // @[pearray.scala 101:13]
  wire [7:0] PE_95_io_data_2_out_bits; // @[pearray.scala 101:13]
  wire  PE_95_io_data_1_in_valid; // @[pearray.scala 101:13]
  wire [7:0] PE_95_io_data_1_in_bits; // @[pearray.scala 101:13]
  wire  PE_95_io_data_1_out_valid; // @[pearray.scala 101:13]
  wire [7:0] PE_95_io_data_1_out_bits; // @[pearray.scala 101:13]
  wire  PE_95_io_data_0_in_valid; // @[pearray.scala 101:13]
  wire [7:0] PE_95_io_data_0_in_bits; // @[pearray.scala 101:13]
  wire  PE_95_io_data_0_out_valid; // @[pearray.scala 101:13]
  wire [7:0] PE_95_io_data_0_out_bits; // @[pearray.scala 101:13]
  wire  PE_95_io_sig_stat2trans; // @[pearray.scala 101:13]
  wire  PE_96_clock; // @[pearray.scala 101:13]
  wire  PE_96_reset; // @[pearray.scala 101:13]
  wire [7:0] PE_96_io_data_2_in_bits; // @[pearray.scala 101:13]
  wire [7:0] PE_96_io_data_2_out_bits; // @[pearray.scala 101:13]
  wire  PE_96_io_data_1_in_valid; // @[pearray.scala 101:13]
  wire [7:0] PE_96_io_data_1_in_bits; // @[pearray.scala 101:13]
  wire  PE_96_io_data_1_out_valid; // @[pearray.scala 101:13]
  wire [7:0] PE_96_io_data_1_out_bits; // @[pearray.scala 101:13]
  wire  PE_96_io_data_0_in_valid; // @[pearray.scala 101:13]
  wire [7:0] PE_96_io_data_0_in_bits; // @[pearray.scala 101:13]
  wire  PE_96_io_data_0_out_valid; // @[pearray.scala 101:13]
  wire [7:0] PE_96_io_data_0_out_bits; // @[pearray.scala 101:13]
  wire  PE_96_io_sig_stat2trans; // @[pearray.scala 101:13]
  wire  PE_97_clock; // @[pearray.scala 101:13]
  wire  PE_97_reset; // @[pearray.scala 101:13]
  wire [7:0] PE_97_io_data_2_in_bits; // @[pearray.scala 101:13]
  wire [7:0] PE_97_io_data_2_out_bits; // @[pearray.scala 101:13]
  wire  PE_97_io_data_1_in_valid; // @[pearray.scala 101:13]
  wire [7:0] PE_97_io_data_1_in_bits; // @[pearray.scala 101:13]
  wire  PE_97_io_data_1_out_valid; // @[pearray.scala 101:13]
  wire [7:0] PE_97_io_data_1_out_bits; // @[pearray.scala 101:13]
  wire  PE_97_io_data_0_in_valid; // @[pearray.scala 101:13]
  wire [7:0] PE_97_io_data_0_in_bits; // @[pearray.scala 101:13]
  wire  PE_97_io_data_0_out_valid; // @[pearray.scala 101:13]
  wire [7:0] PE_97_io_data_0_out_bits; // @[pearray.scala 101:13]
  wire  PE_97_io_sig_stat2trans; // @[pearray.scala 101:13]
  wire  PE_98_clock; // @[pearray.scala 101:13]
  wire  PE_98_reset; // @[pearray.scala 101:13]
  wire [7:0] PE_98_io_data_2_in_bits; // @[pearray.scala 101:13]
  wire [7:0] PE_98_io_data_2_out_bits; // @[pearray.scala 101:13]
  wire  PE_98_io_data_1_in_valid; // @[pearray.scala 101:13]
  wire [7:0] PE_98_io_data_1_in_bits; // @[pearray.scala 101:13]
  wire  PE_98_io_data_1_out_valid; // @[pearray.scala 101:13]
  wire [7:0] PE_98_io_data_1_out_bits; // @[pearray.scala 101:13]
  wire  PE_98_io_data_0_in_valid; // @[pearray.scala 101:13]
  wire [7:0] PE_98_io_data_0_in_bits; // @[pearray.scala 101:13]
  wire  PE_98_io_data_0_out_valid; // @[pearray.scala 101:13]
  wire [7:0] PE_98_io_data_0_out_bits; // @[pearray.scala 101:13]
  wire  PE_98_io_sig_stat2trans; // @[pearray.scala 101:13]
  wire  PE_99_clock; // @[pearray.scala 101:13]
  wire  PE_99_reset; // @[pearray.scala 101:13]
  wire [7:0] PE_99_io_data_2_in_bits; // @[pearray.scala 101:13]
  wire [7:0] PE_99_io_data_2_out_bits; // @[pearray.scala 101:13]
  wire  PE_99_io_data_1_in_valid; // @[pearray.scala 101:13]
  wire [7:0] PE_99_io_data_1_in_bits; // @[pearray.scala 101:13]
  wire  PE_99_io_data_1_out_valid; // @[pearray.scala 101:13]
  wire [7:0] PE_99_io_data_1_out_bits; // @[pearray.scala 101:13]
  wire  PE_99_io_data_0_in_valid; // @[pearray.scala 101:13]
  wire [7:0] PE_99_io_data_0_in_bits; // @[pearray.scala 101:13]
  wire  PE_99_io_data_0_out_valid; // @[pearray.scala 101:13]
  wire [7:0] PE_99_io_data_0_out_bits; // @[pearray.scala 101:13]
  wire  PE_99_io_sig_stat2trans; // @[pearray.scala 101:13]
  wire  PE_100_clock; // @[pearray.scala 101:13]
  wire  PE_100_reset; // @[pearray.scala 101:13]
  wire [7:0] PE_100_io_data_2_in_bits; // @[pearray.scala 101:13]
  wire [7:0] PE_100_io_data_2_out_bits; // @[pearray.scala 101:13]
  wire  PE_100_io_data_1_in_valid; // @[pearray.scala 101:13]
  wire [7:0] PE_100_io_data_1_in_bits; // @[pearray.scala 101:13]
  wire  PE_100_io_data_1_out_valid; // @[pearray.scala 101:13]
  wire [7:0] PE_100_io_data_1_out_bits; // @[pearray.scala 101:13]
  wire  PE_100_io_data_0_in_valid; // @[pearray.scala 101:13]
  wire [7:0] PE_100_io_data_0_in_bits; // @[pearray.scala 101:13]
  wire  PE_100_io_data_0_out_valid; // @[pearray.scala 101:13]
  wire [7:0] PE_100_io_data_0_out_bits; // @[pearray.scala 101:13]
  wire  PE_100_io_sig_stat2trans; // @[pearray.scala 101:13]
  wire  PE_101_clock; // @[pearray.scala 101:13]
  wire  PE_101_reset; // @[pearray.scala 101:13]
  wire [7:0] PE_101_io_data_2_in_bits; // @[pearray.scala 101:13]
  wire [7:0] PE_101_io_data_2_out_bits; // @[pearray.scala 101:13]
  wire  PE_101_io_data_1_in_valid; // @[pearray.scala 101:13]
  wire [7:0] PE_101_io_data_1_in_bits; // @[pearray.scala 101:13]
  wire  PE_101_io_data_1_out_valid; // @[pearray.scala 101:13]
  wire [7:0] PE_101_io_data_1_out_bits; // @[pearray.scala 101:13]
  wire  PE_101_io_data_0_in_valid; // @[pearray.scala 101:13]
  wire [7:0] PE_101_io_data_0_in_bits; // @[pearray.scala 101:13]
  wire  PE_101_io_data_0_out_valid; // @[pearray.scala 101:13]
  wire [7:0] PE_101_io_data_0_out_bits; // @[pearray.scala 101:13]
  wire  PE_101_io_sig_stat2trans; // @[pearray.scala 101:13]
  wire  PE_102_clock; // @[pearray.scala 101:13]
  wire  PE_102_reset; // @[pearray.scala 101:13]
  wire [7:0] PE_102_io_data_2_in_bits; // @[pearray.scala 101:13]
  wire [7:0] PE_102_io_data_2_out_bits; // @[pearray.scala 101:13]
  wire  PE_102_io_data_1_in_valid; // @[pearray.scala 101:13]
  wire [7:0] PE_102_io_data_1_in_bits; // @[pearray.scala 101:13]
  wire  PE_102_io_data_1_out_valid; // @[pearray.scala 101:13]
  wire [7:0] PE_102_io_data_1_out_bits; // @[pearray.scala 101:13]
  wire  PE_102_io_data_0_in_valid; // @[pearray.scala 101:13]
  wire [7:0] PE_102_io_data_0_in_bits; // @[pearray.scala 101:13]
  wire  PE_102_io_data_0_out_valid; // @[pearray.scala 101:13]
  wire [7:0] PE_102_io_data_0_out_bits; // @[pearray.scala 101:13]
  wire  PE_102_io_sig_stat2trans; // @[pearray.scala 101:13]
  wire  PE_103_clock; // @[pearray.scala 101:13]
  wire  PE_103_reset; // @[pearray.scala 101:13]
  wire [7:0] PE_103_io_data_2_in_bits; // @[pearray.scala 101:13]
  wire [7:0] PE_103_io_data_2_out_bits; // @[pearray.scala 101:13]
  wire  PE_103_io_data_1_in_valid; // @[pearray.scala 101:13]
  wire [7:0] PE_103_io_data_1_in_bits; // @[pearray.scala 101:13]
  wire  PE_103_io_data_1_out_valid; // @[pearray.scala 101:13]
  wire [7:0] PE_103_io_data_1_out_bits; // @[pearray.scala 101:13]
  wire  PE_103_io_data_0_in_valid; // @[pearray.scala 101:13]
  wire [7:0] PE_103_io_data_0_in_bits; // @[pearray.scala 101:13]
  wire  PE_103_io_data_0_out_valid; // @[pearray.scala 101:13]
  wire [7:0] PE_103_io_data_0_out_bits; // @[pearray.scala 101:13]
  wire  PE_103_io_sig_stat2trans; // @[pearray.scala 101:13]
  wire  PE_104_clock; // @[pearray.scala 101:13]
  wire  PE_104_reset; // @[pearray.scala 101:13]
  wire [7:0] PE_104_io_data_2_in_bits; // @[pearray.scala 101:13]
  wire [7:0] PE_104_io_data_2_out_bits; // @[pearray.scala 101:13]
  wire  PE_104_io_data_1_in_valid; // @[pearray.scala 101:13]
  wire [7:0] PE_104_io_data_1_in_bits; // @[pearray.scala 101:13]
  wire  PE_104_io_data_1_out_valid; // @[pearray.scala 101:13]
  wire [7:0] PE_104_io_data_1_out_bits; // @[pearray.scala 101:13]
  wire  PE_104_io_data_0_in_valid; // @[pearray.scala 101:13]
  wire [7:0] PE_104_io_data_0_in_bits; // @[pearray.scala 101:13]
  wire  PE_104_io_data_0_out_valid; // @[pearray.scala 101:13]
  wire [7:0] PE_104_io_data_0_out_bits; // @[pearray.scala 101:13]
  wire  PE_104_io_sig_stat2trans; // @[pearray.scala 101:13]
  wire  PE_105_clock; // @[pearray.scala 101:13]
  wire  PE_105_reset; // @[pearray.scala 101:13]
  wire [7:0] PE_105_io_data_2_in_bits; // @[pearray.scala 101:13]
  wire [7:0] PE_105_io_data_2_out_bits; // @[pearray.scala 101:13]
  wire  PE_105_io_data_1_in_valid; // @[pearray.scala 101:13]
  wire [7:0] PE_105_io_data_1_in_bits; // @[pearray.scala 101:13]
  wire  PE_105_io_data_1_out_valid; // @[pearray.scala 101:13]
  wire [7:0] PE_105_io_data_1_out_bits; // @[pearray.scala 101:13]
  wire  PE_105_io_data_0_in_valid; // @[pearray.scala 101:13]
  wire [7:0] PE_105_io_data_0_in_bits; // @[pearray.scala 101:13]
  wire  PE_105_io_data_0_out_valid; // @[pearray.scala 101:13]
  wire [7:0] PE_105_io_data_0_out_bits; // @[pearray.scala 101:13]
  wire  PE_105_io_sig_stat2trans; // @[pearray.scala 101:13]
  wire  PE_106_clock; // @[pearray.scala 101:13]
  wire  PE_106_reset; // @[pearray.scala 101:13]
  wire [7:0] PE_106_io_data_2_in_bits; // @[pearray.scala 101:13]
  wire [7:0] PE_106_io_data_2_out_bits; // @[pearray.scala 101:13]
  wire  PE_106_io_data_1_in_valid; // @[pearray.scala 101:13]
  wire [7:0] PE_106_io_data_1_in_bits; // @[pearray.scala 101:13]
  wire  PE_106_io_data_1_out_valid; // @[pearray.scala 101:13]
  wire [7:0] PE_106_io_data_1_out_bits; // @[pearray.scala 101:13]
  wire  PE_106_io_data_0_in_valid; // @[pearray.scala 101:13]
  wire [7:0] PE_106_io_data_0_in_bits; // @[pearray.scala 101:13]
  wire  PE_106_io_data_0_out_valid; // @[pearray.scala 101:13]
  wire [7:0] PE_106_io_data_0_out_bits; // @[pearray.scala 101:13]
  wire  PE_106_io_sig_stat2trans; // @[pearray.scala 101:13]
  wire  PE_107_clock; // @[pearray.scala 101:13]
  wire  PE_107_reset; // @[pearray.scala 101:13]
  wire [7:0] PE_107_io_data_2_in_bits; // @[pearray.scala 101:13]
  wire [7:0] PE_107_io_data_2_out_bits; // @[pearray.scala 101:13]
  wire  PE_107_io_data_1_in_valid; // @[pearray.scala 101:13]
  wire [7:0] PE_107_io_data_1_in_bits; // @[pearray.scala 101:13]
  wire  PE_107_io_data_1_out_valid; // @[pearray.scala 101:13]
  wire [7:0] PE_107_io_data_1_out_bits; // @[pearray.scala 101:13]
  wire  PE_107_io_data_0_in_valid; // @[pearray.scala 101:13]
  wire [7:0] PE_107_io_data_0_in_bits; // @[pearray.scala 101:13]
  wire  PE_107_io_data_0_out_valid; // @[pearray.scala 101:13]
  wire [7:0] PE_107_io_data_0_out_bits; // @[pearray.scala 101:13]
  wire  PE_107_io_sig_stat2trans; // @[pearray.scala 101:13]
  wire  PE_108_clock; // @[pearray.scala 101:13]
  wire  PE_108_reset; // @[pearray.scala 101:13]
  wire [7:0] PE_108_io_data_2_in_bits; // @[pearray.scala 101:13]
  wire [7:0] PE_108_io_data_2_out_bits; // @[pearray.scala 101:13]
  wire  PE_108_io_data_1_in_valid; // @[pearray.scala 101:13]
  wire [7:0] PE_108_io_data_1_in_bits; // @[pearray.scala 101:13]
  wire  PE_108_io_data_1_out_valid; // @[pearray.scala 101:13]
  wire [7:0] PE_108_io_data_1_out_bits; // @[pearray.scala 101:13]
  wire  PE_108_io_data_0_in_valid; // @[pearray.scala 101:13]
  wire [7:0] PE_108_io_data_0_in_bits; // @[pearray.scala 101:13]
  wire  PE_108_io_data_0_out_valid; // @[pearray.scala 101:13]
  wire [7:0] PE_108_io_data_0_out_bits; // @[pearray.scala 101:13]
  wire  PE_108_io_sig_stat2trans; // @[pearray.scala 101:13]
  wire  PE_109_clock; // @[pearray.scala 101:13]
  wire  PE_109_reset; // @[pearray.scala 101:13]
  wire [7:0] PE_109_io_data_2_in_bits; // @[pearray.scala 101:13]
  wire [7:0] PE_109_io_data_2_out_bits; // @[pearray.scala 101:13]
  wire  PE_109_io_data_1_in_valid; // @[pearray.scala 101:13]
  wire [7:0] PE_109_io_data_1_in_bits; // @[pearray.scala 101:13]
  wire  PE_109_io_data_1_out_valid; // @[pearray.scala 101:13]
  wire [7:0] PE_109_io_data_1_out_bits; // @[pearray.scala 101:13]
  wire  PE_109_io_data_0_in_valid; // @[pearray.scala 101:13]
  wire [7:0] PE_109_io_data_0_in_bits; // @[pearray.scala 101:13]
  wire  PE_109_io_data_0_out_valid; // @[pearray.scala 101:13]
  wire [7:0] PE_109_io_data_0_out_bits; // @[pearray.scala 101:13]
  wire  PE_109_io_sig_stat2trans; // @[pearray.scala 101:13]
  wire  PE_110_clock; // @[pearray.scala 101:13]
  wire  PE_110_reset; // @[pearray.scala 101:13]
  wire [7:0] PE_110_io_data_2_in_bits; // @[pearray.scala 101:13]
  wire [7:0] PE_110_io_data_2_out_bits; // @[pearray.scala 101:13]
  wire  PE_110_io_data_1_in_valid; // @[pearray.scala 101:13]
  wire [7:0] PE_110_io_data_1_in_bits; // @[pearray.scala 101:13]
  wire  PE_110_io_data_1_out_valid; // @[pearray.scala 101:13]
  wire [7:0] PE_110_io_data_1_out_bits; // @[pearray.scala 101:13]
  wire  PE_110_io_data_0_in_valid; // @[pearray.scala 101:13]
  wire [7:0] PE_110_io_data_0_in_bits; // @[pearray.scala 101:13]
  wire  PE_110_io_data_0_out_valid; // @[pearray.scala 101:13]
  wire [7:0] PE_110_io_data_0_out_bits; // @[pearray.scala 101:13]
  wire  PE_110_io_sig_stat2trans; // @[pearray.scala 101:13]
  wire  PE_111_clock; // @[pearray.scala 101:13]
  wire  PE_111_reset; // @[pearray.scala 101:13]
  wire [7:0] PE_111_io_data_2_in_bits; // @[pearray.scala 101:13]
  wire [7:0] PE_111_io_data_2_out_bits; // @[pearray.scala 101:13]
  wire  PE_111_io_data_1_in_valid; // @[pearray.scala 101:13]
  wire [7:0] PE_111_io_data_1_in_bits; // @[pearray.scala 101:13]
  wire  PE_111_io_data_1_out_valid; // @[pearray.scala 101:13]
  wire [7:0] PE_111_io_data_1_out_bits; // @[pearray.scala 101:13]
  wire  PE_111_io_data_0_in_valid; // @[pearray.scala 101:13]
  wire [7:0] PE_111_io_data_0_in_bits; // @[pearray.scala 101:13]
  wire  PE_111_io_data_0_out_valid; // @[pearray.scala 101:13]
  wire [7:0] PE_111_io_data_0_out_bits; // @[pearray.scala 101:13]
  wire  PE_111_io_sig_stat2trans; // @[pearray.scala 101:13]
  wire  PE_112_clock; // @[pearray.scala 101:13]
  wire  PE_112_reset; // @[pearray.scala 101:13]
  wire [7:0] PE_112_io_data_2_in_bits; // @[pearray.scala 101:13]
  wire [7:0] PE_112_io_data_2_out_bits; // @[pearray.scala 101:13]
  wire  PE_112_io_data_1_in_valid; // @[pearray.scala 101:13]
  wire [7:0] PE_112_io_data_1_in_bits; // @[pearray.scala 101:13]
  wire  PE_112_io_data_1_out_valid; // @[pearray.scala 101:13]
  wire [7:0] PE_112_io_data_1_out_bits; // @[pearray.scala 101:13]
  wire  PE_112_io_data_0_in_valid; // @[pearray.scala 101:13]
  wire [7:0] PE_112_io_data_0_in_bits; // @[pearray.scala 101:13]
  wire  PE_112_io_data_0_out_valid; // @[pearray.scala 101:13]
  wire [7:0] PE_112_io_data_0_out_bits; // @[pearray.scala 101:13]
  wire  PE_112_io_sig_stat2trans; // @[pearray.scala 101:13]
  wire  PE_113_clock; // @[pearray.scala 101:13]
  wire  PE_113_reset; // @[pearray.scala 101:13]
  wire [7:0] PE_113_io_data_2_in_bits; // @[pearray.scala 101:13]
  wire [7:0] PE_113_io_data_2_out_bits; // @[pearray.scala 101:13]
  wire  PE_113_io_data_1_in_valid; // @[pearray.scala 101:13]
  wire [7:0] PE_113_io_data_1_in_bits; // @[pearray.scala 101:13]
  wire  PE_113_io_data_1_out_valid; // @[pearray.scala 101:13]
  wire [7:0] PE_113_io_data_1_out_bits; // @[pearray.scala 101:13]
  wire  PE_113_io_data_0_in_valid; // @[pearray.scala 101:13]
  wire [7:0] PE_113_io_data_0_in_bits; // @[pearray.scala 101:13]
  wire  PE_113_io_data_0_out_valid; // @[pearray.scala 101:13]
  wire [7:0] PE_113_io_data_0_out_bits; // @[pearray.scala 101:13]
  wire  PE_113_io_sig_stat2trans; // @[pearray.scala 101:13]
  wire  PE_114_clock; // @[pearray.scala 101:13]
  wire  PE_114_reset; // @[pearray.scala 101:13]
  wire [7:0] PE_114_io_data_2_in_bits; // @[pearray.scala 101:13]
  wire [7:0] PE_114_io_data_2_out_bits; // @[pearray.scala 101:13]
  wire  PE_114_io_data_1_in_valid; // @[pearray.scala 101:13]
  wire [7:0] PE_114_io_data_1_in_bits; // @[pearray.scala 101:13]
  wire  PE_114_io_data_1_out_valid; // @[pearray.scala 101:13]
  wire [7:0] PE_114_io_data_1_out_bits; // @[pearray.scala 101:13]
  wire  PE_114_io_data_0_in_valid; // @[pearray.scala 101:13]
  wire [7:0] PE_114_io_data_0_in_bits; // @[pearray.scala 101:13]
  wire  PE_114_io_data_0_out_valid; // @[pearray.scala 101:13]
  wire [7:0] PE_114_io_data_0_out_bits; // @[pearray.scala 101:13]
  wire  PE_114_io_sig_stat2trans; // @[pearray.scala 101:13]
  wire  PE_115_clock; // @[pearray.scala 101:13]
  wire  PE_115_reset; // @[pearray.scala 101:13]
  wire [7:0] PE_115_io_data_2_in_bits; // @[pearray.scala 101:13]
  wire [7:0] PE_115_io_data_2_out_bits; // @[pearray.scala 101:13]
  wire  PE_115_io_data_1_in_valid; // @[pearray.scala 101:13]
  wire [7:0] PE_115_io_data_1_in_bits; // @[pearray.scala 101:13]
  wire  PE_115_io_data_1_out_valid; // @[pearray.scala 101:13]
  wire [7:0] PE_115_io_data_1_out_bits; // @[pearray.scala 101:13]
  wire  PE_115_io_data_0_in_valid; // @[pearray.scala 101:13]
  wire [7:0] PE_115_io_data_0_in_bits; // @[pearray.scala 101:13]
  wire  PE_115_io_data_0_out_valid; // @[pearray.scala 101:13]
  wire [7:0] PE_115_io_data_0_out_bits; // @[pearray.scala 101:13]
  wire  PE_115_io_sig_stat2trans; // @[pearray.scala 101:13]
  wire  PE_116_clock; // @[pearray.scala 101:13]
  wire  PE_116_reset; // @[pearray.scala 101:13]
  wire [7:0] PE_116_io_data_2_in_bits; // @[pearray.scala 101:13]
  wire [7:0] PE_116_io_data_2_out_bits; // @[pearray.scala 101:13]
  wire  PE_116_io_data_1_in_valid; // @[pearray.scala 101:13]
  wire [7:0] PE_116_io_data_1_in_bits; // @[pearray.scala 101:13]
  wire  PE_116_io_data_1_out_valid; // @[pearray.scala 101:13]
  wire [7:0] PE_116_io_data_1_out_bits; // @[pearray.scala 101:13]
  wire  PE_116_io_data_0_in_valid; // @[pearray.scala 101:13]
  wire [7:0] PE_116_io_data_0_in_bits; // @[pearray.scala 101:13]
  wire  PE_116_io_data_0_out_valid; // @[pearray.scala 101:13]
  wire [7:0] PE_116_io_data_0_out_bits; // @[pearray.scala 101:13]
  wire  PE_116_io_sig_stat2trans; // @[pearray.scala 101:13]
  wire  PE_117_clock; // @[pearray.scala 101:13]
  wire  PE_117_reset; // @[pearray.scala 101:13]
  wire [7:0] PE_117_io_data_2_in_bits; // @[pearray.scala 101:13]
  wire [7:0] PE_117_io_data_2_out_bits; // @[pearray.scala 101:13]
  wire  PE_117_io_data_1_in_valid; // @[pearray.scala 101:13]
  wire [7:0] PE_117_io_data_1_in_bits; // @[pearray.scala 101:13]
  wire  PE_117_io_data_1_out_valid; // @[pearray.scala 101:13]
  wire [7:0] PE_117_io_data_1_out_bits; // @[pearray.scala 101:13]
  wire  PE_117_io_data_0_in_valid; // @[pearray.scala 101:13]
  wire [7:0] PE_117_io_data_0_in_bits; // @[pearray.scala 101:13]
  wire  PE_117_io_data_0_out_valid; // @[pearray.scala 101:13]
  wire [7:0] PE_117_io_data_0_out_bits; // @[pearray.scala 101:13]
  wire  PE_117_io_sig_stat2trans; // @[pearray.scala 101:13]
  wire  PE_118_clock; // @[pearray.scala 101:13]
  wire  PE_118_reset; // @[pearray.scala 101:13]
  wire [7:0] PE_118_io_data_2_in_bits; // @[pearray.scala 101:13]
  wire [7:0] PE_118_io_data_2_out_bits; // @[pearray.scala 101:13]
  wire  PE_118_io_data_1_in_valid; // @[pearray.scala 101:13]
  wire [7:0] PE_118_io_data_1_in_bits; // @[pearray.scala 101:13]
  wire  PE_118_io_data_1_out_valid; // @[pearray.scala 101:13]
  wire [7:0] PE_118_io_data_1_out_bits; // @[pearray.scala 101:13]
  wire  PE_118_io_data_0_in_valid; // @[pearray.scala 101:13]
  wire [7:0] PE_118_io_data_0_in_bits; // @[pearray.scala 101:13]
  wire  PE_118_io_data_0_out_valid; // @[pearray.scala 101:13]
  wire [7:0] PE_118_io_data_0_out_bits; // @[pearray.scala 101:13]
  wire  PE_118_io_sig_stat2trans; // @[pearray.scala 101:13]
  wire  PE_119_clock; // @[pearray.scala 101:13]
  wire  PE_119_reset; // @[pearray.scala 101:13]
  wire [7:0] PE_119_io_data_2_in_bits; // @[pearray.scala 101:13]
  wire [7:0] PE_119_io_data_2_out_bits; // @[pearray.scala 101:13]
  wire  PE_119_io_data_1_in_valid; // @[pearray.scala 101:13]
  wire [7:0] PE_119_io_data_1_in_bits; // @[pearray.scala 101:13]
  wire  PE_119_io_data_1_out_valid; // @[pearray.scala 101:13]
  wire [7:0] PE_119_io_data_1_out_bits; // @[pearray.scala 101:13]
  wire  PE_119_io_data_0_in_valid; // @[pearray.scala 101:13]
  wire [7:0] PE_119_io_data_0_in_bits; // @[pearray.scala 101:13]
  wire  PE_119_io_data_0_out_valid; // @[pearray.scala 101:13]
  wire [7:0] PE_119_io_data_0_out_bits; // @[pearray.scala 101:13]
  wire  PE_119_io_sig_stat2trans; // @[pearray.scala 101:13]
  wire  PE_120_clock; // @[pearray.scala 101:13]
  wire  PE_120_reset; // @[pearray.scala 101:13]
  wire [7:0] PE_120_io_data_2_in_bits; // @[pearray.scala 101:13]
  wire [7:0] PE_120_io_data_2_out_bits; // @[pearray.scala 101:13]
  wire  PE_120_io_data_1_in_valid; // @[pearray.scala 101:13]
  wire [7:0] PE_120_io_data_1_in_bits; // @[pearray.scala 101:13]
  wire  PE_120_io_data_1_out_valid; // @[pearray.scala 101:13]
  wire [7:0] PE_120_io_data_1_out_bits; // @[pearray.scala 101:13]
  wire  PE_120_io_data_0_in_valid; // @[pearray.scala 101:13]
  wire [7:0] PE_120_io_data_0_in_bits; // @[pearray.scala 101:13]
  wire  PE_120_io_data_0_out_valid; // @[pearray.scala 101:13]
  wire [7:0] PE_120_io_data_0_out_bits; // @[pearray.scala 101:13]
  wire  PE_120_io_sig_stat2trans; // @[pearray.scala 101:13]
  wire  PE_121_clock; // @[pearray.scala 101:13]
  wire  PE_121_reset; // @[pearray.scala 101:13]
  wire [7:0] PE_121_io_data_2_in_bits; // @[pearray.scala 101:13]
  wire [7:0] PE_121_io_data_2_out_bits; // @[pearray.scala 101:13]
  wire  PE_121_io_data_1_in_valid; // @[pearray.scala 101:13]
  wire [7:0] PE_121_io_data_1_in_bits; // @[pearray.scala 101:13]
  wire  PE_121_io_data_1_out_valid; // @[pearray.scala 101:13]
  wire [7:0] PE_121_io_data_1_out_bits; // @[pearray.scala 101:13]
  wire  PE_121_io_data_0_in_valid; // @[pearray.scala 101:13]
  wire [7:0] PE_121_io_data_0_in_bits; // @[pearray.scala 101:13]
  wire  PE_121_io_data_0_out_valid; // @[pearray.scala 101:13]
  wire [7:0] PE_121_io_data_0_out_bits; // @[pearray.scala 101:13]
  wire  PE_121_io_sig_stat2trans; // @[pearray.scala 101:13]
  wire  PE_122_clock; // @[pearray.scala 101:13]
  wire  PE_122_reset; // @[pearray.scala 101:13]
  wire [7:0] PE_122_io_data_2_in_bits; // @[pearray.scala 101:13]
  wire [7:0] PE_122_io_data_2_out_bits; // @[pearray.scala 101:13]
  wire  PE_122_io_data_1_in_valid; // @[pearray.scala 101:13]
  wire [7:0] PE_122_io_data_1_in_bits; // @[pearray.scala 101:13]
  wire  PE_122_io_data_1_out_valid; // @[pearray.scala 101:13]
  wire [7:0] PE_122_io_data_1_out_bits; // @[pearray.scala 101:13]
  wire  PE_122_io_data_0_in_valid; // @[pearray.scala 101:13]
  wire [7:0] PE_122_io_data_0_in_bits; // @[pearray.scala 101:13]
  wire  PE_122_io_data_0_out_valid; // @[pearray.scala 101:13]
  wire [7:0] PE_122_io_data_0_out_bits; // @[pearray.scala 101:13]
  wire  PE_122_io_sig_stat2trans; // @[pearray.scala 101:13]
  wire  PE_123_clock; // @[pearray.scala 101:13]
  wire  PE_123_reset; // @[pearray.scala 101:13]
  wire [7:0] PE_123_io_data_2_in_bits; // @[pearray.scala 101:13]
  wire [7:0] PE_123_io_data_2_out_bits; // @[pearray.scala 101:13]
  wire  PE_123_io_data_1_in_valid; // @[pearray.scala 101:13]
  wire [7:0] PE_123_io_data_1_in_bits; // @[pearray.scala 101:13]
  wire  PE_123_io_data_1_out_valid; // @[pearray.scala 101:13]
  wire [7:0] PE_123_io_data_1_out_bits; // @[pearray.scala 101:13]
  wire  PE_123_io_data_0_in_valid; // @[pearray.scala 101:13]
  wire [7:0] PE_123_io_data_0_in_bits; // @[pearray.scala 101:13]
  wire  PE_123_io_data_0_out_valid; // @[pearray.scala 101:13]
  wire [7:0] PE_123_io_data_0_out_bits; // @[pearray.scala 101:13]
  wire  PE_123_io_sig_stat2trans; // @[pearray.scala 101:13]
  wire  PE_124_clock; // @[pearray.scala 101:13]
  wire  PE_124_reset; // @[pearray.scala 101:13]
  wire [7:0] PE_124_io_data_2_in_bits; // @[pearray.scala 101:13]
  wire [7:0] PE_124_io_data_2_out_bits; // @[pearray.scala 101:13]
  wire  PE_124_io_data_1_in_valid; // @[pearray.scala 101:13]
  wire [7:0] PE_124_io_data_1_in_bits; // @[pearray.scala 101:13]
  wire  PE_124_io_data_1_out_valid; // @[pearray.scala 101:13]
  wire [7:0] PE_124_io_data_1_out_bits; // @[pearray.scala 101:13]
  wire  PE_124_io_data_0_in_valid; // @[pearray.scala 101:13]
  wire [7:0] PE_124_io_data_0_in_bits; // @[pearray.scala 101:13]
  wire  PE_124_io_data_0_out_valid; // @[pearray.scala 101:13]
  wire [7:0] PE_124_io_data_0_out_bits; // @[pearray.scala 101:13]
  wire  PE_124_io_sig_stat2trans; // @[pearray.scala 101:13]
  wire  PE_125_clock; // @[pearray.scala 101:13]
  wire  PE_125_reset; // @[pearray.scala 101:13]
  wire [7:0] PE_125_io_data_2_in_bits; // @[pearray.scala 101:13]
  wire [7:0] PE_125_io_data_2_out_bits; // @[pearray.scala 101:13]
  wire  PE_125_io_data_1_in_valid; // @[pearray.scala 101:13]
  wire [7:0] PE_125_io_data_1_in_bits; // @[pearray.scala 101:13]
  wire  PE_125_io_data_1_out_valid; // @[pearray.scala 101:13]
  wire [7:0] PE_125_io_data_1_out_bits; // @[pearray.scala 101:13]
  wire  PE_125_io_data_0_in_valid; // @[pearray.scala 101:13]
  wire [7:0] PE_125_io_data_0_in_bits; // @[pearray.scala 101:13]
  wire  PE_125_io_data_0_out_valid; // @[pearray.scala 101:13]
  wire [7:0] PE_125_io_data_0_out_bits; // @[pearray.scala 101:13]
  wire  PE_125_io_sig_stat2trans; // @[pearray.scala 101:13]
  wire  PE_126_clock; // @[pearray.scala 101:13]
  wire  PE_126_reset; // @[pearray.scala 101:13]
  wire [7:0] PE_126_io_data_2_in_bits; // @[pearray.scala 101:13]
  wire [7:0] PE_126_io_data_2_out_bits; // @[pearray.scala 101:13]
  wire  PE_126_io_data_1_in_valid; // @[pearray.scala 101:13]
  wire [7:0] PE_126_io_data_1_in_bits; // @[pearray.scala 101:13]
  wire  PE_126_io_data_1_out_valid; // @[pearray.scala 101:13]
  wire [7:0] PE_126_io_data_1_out_bits; // @[pearray.scala 101:13]
  wire  PE_126_io_data_0_in_valid; // @[pearray.scala 101:13]
  wire [7:0] PE_126_io_data_0_in_bits; // @[pearray.scala 101:13]
  wire  PE_126_io_data_0_out_valid; // @[pearray.scala 101:13]
  wire [7:0] PE_126_io_data_0_out_bits; // @[pearray.scala 101:13]
  wire  PE_126_io_sig_stat2trans; // @[pearray.scala 101:13]
  wire  PE_127_clock; // @[pearray.scala 101:13]
  wire  PE_127_reset; // @[pearray.scala 101:13]
  wire [7:0] PE_127_io_data_2_in_bits; // @[pearray.scala 101:13]
  wire [7:0] PE_127_io_data_2_out_bits; // @[pearray.scala 101:13]
  wire  PE_127_io_data_1_in_valid; // @[pearray.scala 101:13]
  wire [7:0] PE_127_io_data_1_in_bits; // @[pearray.scala 101:13]
  wire  PE_127_io_data_1_out_valid; // @[pearray.scala 101:13]
  wire [7:0] PE_127_io_data_1_out_bits; // @[pearray.scala 101:13]
  wire  PE_127_io_data_0_in_valid; // @[pearray.scala 101:13]
  wire [7:0] PE_127_io_data_0_in_bits; // @[pearray.scala 101:13]
  wire  PE_127_io_data_0_out_valid; // @[pearray.scala 101:13]
  wire [7:0] PE_127_io_data_0_out_bits; // @[pearray.scala 101:13]
  wire  PE_127_io_sig_stat2trans; // @[pearray.scala 101:13]
  wire  PENetwork_io_to_pes_0_out_valid; // @[pearray.scala 134:13]
  wire [7:0] PENetwork_io_to_pes_0_out_bits; // @[pearray.scala 134:13]
  wire  PENetwork_io_to_pes_1_in_valid; // @[pearray.scala 134:13]
  wire [7:0] PENetwork_io_to_pes_1_in_bits; // @[pearray.scala 134:13]
  wire  PENetwork_io_to_pes_1_out_valid; // @[pearray.scala 134:13]
  wire [7:0] PENetwork_io_to_pes_1_out_bits; // @[pearray.scala 134:13]
  wire  PENetwork_io_to_pes_2_in_valid; // @[pearray.scala 134:13]
  wire [7:0] PENetwork_io_to_pes_2_in_bits; // @[pearray.scala 134:13]
  wire  PENetwork_io_to_pes_2_out_valid; // @[pearray.scala 134:13]
  wire [7:0] PENetwork_io_to_pes_2_out_bits; // @[pearray.scala 134:13]
  wire  PENetwork_io_to_pes_3_in_valid; // @[pearray.scala 134:13]
  wire [7:0] PENetwork_io_to_pes_3_in_bits; // @[pearray.scala 134:13]
  wire  PENetwork_io_to_pes_3_out_valid; // @[pearray.scala 134:13]
  wire [7:0] PENetwork_io_to_pes_3_out_bits; // @[pearray.scala 134:13]
  wire  PENetwork_io_to_pes_4_in_valid; // @[pearray.scala 134:13]
  wire [7:0] PENetwork_io_to_pes_4_in_bits; // @[pearray.scala 134:13]
  wire  PENetwork_io_to_pes_4_out_valid; // @[pearray.scala 134:13]
  wire [7:0] PENetwork_io_to_pes_4_out_bits; // @[pearray.scala 134:13]
  wire  PENetwork_io_to_pes_5_in_valid; // @[pearray.scala 134:13]
  wire [7:0] PENetwork_io_to_pes_5_in_bits; // @[pearray.scala 134:13]
  wire  PENetwork_io_to_pes_5_out_valid; // @[pearray.scala 134:13]
  wire [7:0] PENetwork_io_to_pes_5_out_bits; // @[pearray.scala 134:13]
  wire  PENetwork_io_to_pes_6_in_valid; // @[pearray.scala 134:13]
  wire [7:0] PENetwork_io_to_pes_6_in_bits; // @[pearray.scala 134:13]
  wire  PENetwork_io_to_pes_6_out_valid; // @[pearray.scala 134:13]
  wire [7:0] PENetwork_io_to_pes_6_out_bits; // @[pearray.scala 134:13]
  wire  PENetwork_io_to_pes_7_in_valid; // @[pearray.scala 134:13]
  wire [7:0] PENetwork_io_to_pes_7_in_bits; // @[pearray.scala 134:13]
  wire  PENetwork_io_to_pes_7_out_valid; // @[pearray.scala 134:13]
  wire [7:0] PENetwork_io_to_pes_7_out_bits; // @[pearray.scala 134:13]
  wire  PENetwork_io_to_mem_valid; // @[pearray.scala 134:13]
  wire [7:0] PENetwork_io_to_mem_bits; // @[pearray.scala 134:13]
  wire  PENetwork_1_io_to_pes_0_out_valid; // @[pearray.scala 134:13]
  wire [7:0] PENetwork_1_io_to_pes_0_out_bits; // @[pearray.scala 134:13]
  wire  PENetwork_1_io_to_pes_1_in_valid; // @[pearray.scala 134:13]
  wire [7:0] PENetwork_1_io_to_pes_1_in_bits; // @[pearray.scala 134:13]
  wire  PENetwork_1_io_to_pes_1_out_valid; // @[pearray.scala 134:13]
  wire [7:0] PENetwork_1_io_to_pes_1_out_bits; // @[pearray.scala 134:13]
  wire  PENetwork_1_io_to_pes_2_in_valid; // @[pearray.scala 134:13]
  wire [7:0] PENetwork_1_io_to_pes_2_in_bits; // @[pearray.scala 134:13]
  wire  PENetwork_1_io_to_pes_2_out_valid; // @[pearray.scala 134:13]
  wire [7:0] PENetwork_1_io_to_pes_2_out_bits; // @[pearray.scala 134:13]
  wire  PENetwork_1_io_to_pes_3_in_valid; // @[pearray.scala 134:13]
  wire [7:0] PENetwork_1_io_to_pes_3_in_bits; // @[pearray.scala 134:13]
  wire  PENetwork_1_io_to_pes_3_out_valid; // @[pearray.scala 134:13]
  wire [7:0] PENetwork_1_io_to_pes_3_out_bits; // @[pearray.scala 134:13]
  wire  PENetwork_1_io_to_pes_4_in_valid; // @[pearray.scala 134:13]
  wire [7:0] PENetwork_1_io_to_pes_4_in_bits; // @[pearray.scala 134:13]
  wire  PENetwork_1_io_to_pes_4_out_valid; // @[pearray.scala 134:13]
  wire [7:0] PENetwork_1_io_to_pes_4_out_bits; // @[pearray.scala 134:13]
  wire  PENetwork_1_io_to_pes_5_in_valid; // @[pearray.scala 134:13]
  wire [7:0] PENetwork_1_io_to_pes_5_in_bits; // @[pearray.scala 134:13]
  wire  PENetwork_1_io_to_pes_5_out_valid; // @[pearray.scala 134:13]
  wire [7:0] PENetwork_1_io_to_pes_5_out_bits; // @[pearray.scala 134:13]
  wire  PENetwork_1_io_to_pes_6_in_valid; // @[pearray.scala 134:13]
  wire [7:0] PENetwork_1_io_to_pes_6_in_bits; // @[pearray.scala 134:13]
  wire  PENetwork_1_io_to_pes_6_out_valid; // @[pearray.scala 134:13]
  wire [7:0] PENetwork_1_io_to_pes_6_out_bits; // @[pearray.scala 134:13]
  wire  PENetwork_1_io_to_pes_7_in_valid; // @[pearray.scala 134:13]
  wire [7:0] PENetwork_1_io_to_pes_7_in_bits; // @[pearray.scala 134:13]
  wire  PENetwork_1_io_to_pes_7_out_valid; // @[pearray.scala 134:13]
  wire [7:0] PENetwork_1_io_to_pes_7_out_bits; // @[pearray.scala 134:13]
  wire  PENetwork_1_io_to_mem_valid; // @[pearray.scala 134:13]
  wire [7:0] PENetwork_1_io_to_mem_bits; // @[pearray.scala 134:13]
  wire  PENetwork_2_io_to_pes_0_out_valid; // @[pearray.scala 134:13]
  wire [7:0] PENetwork_2_io_to_pes_0_out_bits; // @[pearray.scala 134:13]
  wire  PENetwork_2_io_to_pes_1_in_valid; // @[pearray.scala 134:13]
  wire [7:0] PENetwork_2_io_to_pes_1_in_bits; // @[pearray.scala 134:13]
  wire  PENetwork_2_io_to_pes_1_out_valid; // @[pearray.scala 134:13]
  wire [7:0] PENetwork_2_io_to_pes_1_out_bits; // @[pearray.scala 134:13]
  wire  PENetwork_2_io_to_pes_2_in_valid; // @[pearray.scala 134:13]
  wire [7:0] PENetwork_2_io_to_pes_2_in_bits; // @[pearray.scala 134:13]
  wire  PENetwork_2_io_to_pes_2_out_valid; // @[pearray.scala 134:13]
  wire [7:0] PENetwork_2_io_to_pes_2_out_bits; // @[pearray.scala 134:13]
  wire  PENetwork_2_io_to_pes_3_in_valid; // @[pearray.scala 134:13]
  wire [7:0] PENetwork_2_io_to_pes_3_in_bits; // @[pearray.scala 134:13]
  wire  PENetwork_2_io_to_pes_3_out_valid; // @[pearray.scala 134:13]
  wire [7:0] PENetwork_2_io_to_pes_3_out_bits; // @[pearray.scala 134:13]
  wire  PENetwork_2_io_to_pes_4_in_valid; // @[pearray.scala 134:13]
  wire [7:0] PENetwork_2_io_to_pes_4_in_bits; // @[pearray.scala 134:13]
  wire  PENetwork_2_io_to_pes_4_out_valid; // @[pearray.scala 134:13]
  wire [7:0] PENetwork_2_io_to_pes_4_out_bits; // @[pearray.scala 134:13]
  wire  PENetwork_2_io_to_pes_5_in_valid; // @[pearray.scala 134:13]
  wire [7:0] PENetwork_2_io_to_pes_5_in_bits; // @[pearray.scala 134:13]
  wire  PENetwork_2_io_to_pes_5_out_valid; // @[pearray.scala 134:13]
  wire [7:0] PENetwork_2_io_to_pes_5_out_bits; // @[pearray.scala 134:13]
  wire  PENetwork_2_io_to_pes_6_in_valid; // @[pearray.scala 134:13]
  wire [7:0] PENetwork_2_io_to_pes_6_in_bits; // @[pearray.scala 134:13]
  wire  PENetwork_2_io_to_pes_6_out_valid; // @[pearray.scala 134:13]
  wire [7:0] PENetwork_2_io_to_pes_6_out_bits; // @[pearray.scala 134:13]
  wire  PENetwork_2_io_to_pes_7_in_valid; // @[pearray.scala 134:13]
  wire [7:0] PENetwork_2_io_to_pes_7_in_bits; // @[pearray.scala 134:13]
  wire  PENetwork_2_io_to_pes_7_out_valid; // @[pearray.scala 134:13]
  wire [7:0] PENetwork_2_io_to_pes_7_out_bits; // @[pearray.scala 134:13]
  wire  PENetwork_2_io_to_mem_valid; // @[pearray.scala 134:13]
  wire [7:0] PENetwork_2_io_to_mem_bits; // @[pearray.scala 134:13]
  wire  PENetwork_3_io_to_pes_0_out_valid; // @[pearray.scala 134:13]
  wire [7:0] PENetwork_3_io_to_pes_0_out_bits; // @[pearray.scala 134:13]
  wire  PENetwork_3_io_to_pes_1_in_valid; // @[pearray.scala 134:13]
  wire [7:0] PENetwork_3_io_to_pes_1_in_bits; // @[pearray.scala 134:13]
  wire  PENetwork_3_io_to_pes_1_out_valid; // @[pearray.scala 134:13]
  wire [7:0] PENetwork_3_io_to_pes_1_out_bits; // @[pearray.scala 134:13]
  wire  PENetwork_3_io_to_pes_2_in_valid; // @[pearray.scala 134:13]
  wire [7:0] PENetwork_3_io_to_pes_2_in_bits; // @[pearray.scala 134:13]
  wire  PENetwork_3_io_to_pes_2_out_valid; // @[pearray.scala 134:13]
  wire [7:0] PENetwork_3_io_to_pes_2_out_bits; // @[pearray.scala 134:13]
  wire  PENetwork_3_io_to_pes_3_in_valid; // @[pearray.scala 134:13]
  wire [7:0] PENetwork_3_io_to_pes_3_in_bits; // @[pearray.scala 134:13]
  wire  PENetwork_3_io_to_pes_3_out_valid; // @[pearray.scala 134:13]
  wire [7:0] PENetwork_3_io_to_pes_3_out_bits; // @[pearray.scala 134:13]
  wire  PENetwork_3_io_to_pes_4_in_valid; // @[pearray.scala 134:13]
  wire [7:0] PENetwork_3_io_to_pes_4_in_bits; // @[pearray.scala 134:13]
  wire  PENetwork_3_io_to_pes_4_out_valid; // @[pearray.scala 134:13]
  wire [7:0] PENetwork_3_io_to_pes_4_out_bits; // @[pearray.scala 134:13]
  wire  PENetwork_3_io_to_pes_5_in_valid; // @[pearray.scala 134:13]
  wire [7:0] PENetwork_3_io_to_pes_5_in_bits; // @[pearray.scala 134:13]
  wire  PENetwork_3_io_to_pes_5_out_valid; // @[pearray.scala 134:13]
  wire [7:0] PENetwork_3_io_to_pes_5_out_bits; // @[pearray.scala 134:13]
  wire  PENetwork_3_io_to_pes_6_in_valid; // @[pearray.scala 134:13]
  wire [7:0] PENetwork_3_io_to_pes_6_in_bits; // @[pearray.scala 134:13]
  wire  PENetwork_3_io_to_pes_6_out_valid; // @[pearray.scala 134:13]
  wire [7:0] PENetwork_3_io_to_pes_6_out_bits; // @[pearray.scala 134:13]
  wire  PENetwork_3_io_to_pes_7_in_valid; // @[pearray.scala 134:13]
  wire [7:0] PENetwork_3_io_to_pes_7_in_bits; // @[pearray.scala 134:13]
  wire  PENetwork_3_io_to_pes_7_out_valid; // @[pearray.scala 134:13]
  wire [7:0] PENetwork_3_io_to_pes_7_out_bits; // @[pearray.scala 134:13]
  wire  PENetwork_3_io_to_mem_valid; // @[pearray.scala 134:13]
  wire [7:0] PENetwork_3_io_to_mem_bits; // @[pearray.scala 134:13]
  wire  PENetwork_4_io_to_pes_0_out_valid; // @[pearray.scala 134:13]
  wire [7:0] PENetwork_4_io_to_pes_0_out_bits; // @[pearray.scala 134:13]
  wire  PENetwork_4_io_to_pes_1_in_valid; // @[pearray.scala 134:13]
  wire [7:0] PENetwork_4_io_to_pes_1_in_bits; // @[pearray.scala 134:13]
  wire  PENetwork_4_io_to_pes_1_out_valid; // @[pearray.scala 134:13]
  wire [7:0] PENetwork_4_io_to_pes_1_out_bits; // @[pearray.scala 134:13]
  wire  PENetwork_4_io_to_pes_2_in_valid; // @[pearray.scala 134:13]
  wire [7:0] PENetwork_4_io_to_pes_2_in_bits; // @[pearray.scala 134:13]
  wire  PENetwork_4_io_to_pes_2_out_valid; // @[pearray.scala 134:13]
  wire [7:0] PENetwork_4_io_to_pes_2_out_bits; // @[pearray.scala 134:13]
  wire  PENetwork_4_io_to_pes_3_in_valid; // @[pearray.scala 134:13]
  wire [7:0] PENetwork_4_io_to_pes_3_in_bits; // @[pearray.scala 134:13]
  wire  PENetwork_4_io_to_pes_3_out_valid; // @[pearray.scala 134:13]
  wire [7:0] PENetwork_4_io_to_pes_3_out_bits; // @[pearray.scala 134:13]
  wire  PENetwork_4_io_to_pes_4_in_valid; // @[pearray.scala 134:13]
  wire [7:0] PENetwork_4_io_to_pes_4_in_bits; // @[pearray.scala 134:13]
  wire  PENetwork_4_io_to_pes_4_out_valid; // @[pearray.scala 134:13]
  wire [7:0] PENetwork_4_io_to_pes_4_out_bits; // @[pearray.scala 134:13]
  wire  PENetwork_4_io_to_pes_5_in_valid; // @[pearray.scala 134:13]
  wire [7:0] PENetwork_4_io_to_pes_5_in_bits; // @[pearray.scala 134:13]
  wire  PENetwork_4_io_to_pes_5_out_valid; // @[pearray.scala 134:13]
  wire [7:0] PENetwork_4_io_to_pes_5_out_bits; // @[pearray.scala 134:13]
  wire  PENetwork_4_io_to_pes_6_in_valid; // @[pearray.scala 134:13]
  wire [7:0] PENetwork_4_io_to_pes_6_in_bits; // @[pearray.scala 134:13]
  wire  PENetwork_4_io_to_pes_6_out_valid; // @[pearray.scala 134:13]
  wire [7:0] PENetwork_4_io_to_pes_6_out_bits; // @[pearray.scala 134:13]
  wire  PENetwork_4_io_to_pes_7_in_valid; // @[pearray.scala 134:13]
  wire [7:0] PENetwork_4_io_to_pes_7_in_bits; // @[pearray.scala 134:13]
  wire  PENetwork_4_io_to_pes_7_out_valid; // @[pearray.scala 134:13]
  wire [7:0] PENetwork_4_io_to_pes_7_out_bits; // @[pearray.scala 134:13]
  wire  PENetwork_4_io_to_mem_valid; // @[pearray.scala 134:13]
  wire [7:0] PENetwork_4_io_to_mem_bits; // @[pearray.scala 134:13]
  wire  PENetwork_5_io_to_pes_0_out_valid; // @[pearray.scala 134:13]
  wire [7:0] PENetwork_5_io_to_pes_0_out_bits; // @[pearray.scala 134:13]
  wire  PENetwork_5_io_to_pes_1_in_valid; // @[pearray.scala 134:13]
  wire [7:0] PENetwork_5_io_to_pes_1_in_bits; // @[pearray.scala 134:13]
  wire  PENetwork_5_io_to_pes_1_out_valid; // @[pearray.scala 134:13]
  wire [7:0] PENetwork_5_io_to_pes_1_out_bits; // @[pearray.scala 134:13]
  wire  PENetwork_5_io_to_pes_2_in_valid; // @[pearray.scala 134:13]
  wire [7:0] PENetwork_5_io_to_pes_2_in_bits; // @[pearray.scala 134:13]
  wire  PENetwork_5_io_to_pes_2_out_valid; // @[pearray.scala 134:13]
  wire [7:0] PENetwork_5_io_to_pes_2_out_bits; // @[pearray.scala 134:13]
  wire  PENetwork_5_io_to_pes_3_in_valid; // @[pearray.scala 134:13]
  wire [7:0] PENetwork_5_io_to_pes_3_in_bits; // @[pearray.scala 134:13]
  wire  PENetwork_5_io_to_pes_3_out_valid; // @[pearray.scala 134:13]
  wire [7:0] PENetwork_5_io_to_pes_3_out_bits; // @[pearray.scala 134:13]
  wire  PENetwork_5_io_to_pes_4_in_valid; // @[pearray.scala 134:13]
  wire [7:0] PENetwork_5_io_to_pes_4_in_bits; // @[pearray.scala 134:13]
  wire  PENetwork_5_io_to_pes_4_out_valid; // @[pearray.scala 134:13]
  wire [7:0] PENetwork_5_io_to_pes_4_out_bits; // @[pearray.scala 134:13]
  wire  PENetwork_5_io_to_pes_5_in_valid; // @[pearray.scala 134:13]
  wire [7:0] PENetwork_5_io_to_pes_5_in_bits; // @[pearray.scala 134:13]
  wire  PENetwork_5_io_to_pes_5_out_valid; // @[pearray.scala 134:13]
  wire [7:0] PENetwork_5_io_to_pes_5_out_bits; // @[pearray.scala 134:13]
  wire  PENetwork_5_io_to_pes_6_in_valid; // @[pearray.scala 134:13]
  wire [7:0] PENetwork_5_io_to_pes_6_in_bits; // @[pearray.scala 134:13]
  wire  PENetwork_5_io_to_pes_6_out_valid; // @[pearray.scala 134:13]
  wire [7:0] PENetwork_5_io_to_pes_6_out_bits; // @[pearray.scala 134:13]
  wire  PENetwork_5_io_to_pes_7_in_valid; // @[pearray.scala 134:13]
  wire [7:0] PENetwork_5_io_to_pes_7_in_bits; // @[pearray.scala 134:13]
  wire  PENetwork_5_io_to_pes_7_out_valid; // @[pearray.scala 134:13]
  wire [7:0] PENetwork_5_io_to_pes_7_out_bits; // @[pearray.scala 134:13]
  wire  PENetwork_5_io_to_mem_valid; // @[pearray.scala 134:13]
  wire [7:0] PENetwork_5_io_to_mem_bits; // @[pearray.scala 134:13]
  wire  PENetwork_6_io_to_pes_0_out_valid; // @[pearray.scala 134:13]
  wire [7:0] PENetwork_6_io_to_pes_0_out_bits; // @[pearray.scala 134:13]
  wire  PENetwork_6_io_to_pes_1_in_valid; // @[pearray.scala 134:13]
  wire [7:0] PENetwork_6_io_to_pes_1_in_bits; // @[pearray.scala 134:13]
  wire  PENetwork_6_io_to_pes_1_out_valid; // @[pearray.scala 134:13]
  wire [7:0] PENetwork_6_io_to_pes_1_out_bits; // @[pearray.scala 134:13]
  wire  PENetwork_6_io_to_pes_2_in_valid; // @[pearray.scala 134:13]
  wire [7:0] PENetwork_6_io_to_pes_2_in_bits; // @[pearray.scala 134:13]
  wire  PENetwork_6_io_to_pes_2_out_valid; // @[pearray.scala 134:13]
  wire [7:0] PENetwork_6_io_to_pes_2_out_bits; // @[pearray.scala 134:13]
  wire  PENetwork_6_io_to_pes_3_in_valid; // @[pearray.scala 134:13]
  wire [7:0] PENetwork_6_io_to_pes_3_in_bits; // @[pearray.scala 134:13]
  wire  PENetwork_6_io_to_pes_3_out_valid; // @[pearray.scala 134:13]
  wire [7:0] PENetwork_6_io_to_pes_3_out_bits; // @[pearray.scala 134:13]
  wire  PENetwork_6_io_to_pes_4_in_valid; // @[pearray.scala 134:13]
  wire [7:0] PENetwork_6_io_to_pes_4_in_bits; // @[pearray.scala 134:13]
  wire  PENetwork_6_io_to_pes_4_out_valid; // @[pearray.scala 134:13]
  wire [7:0] PENetwork_6_io_to_pes_4_out_bits; // @[pearray.scala 134:13]
  wire  PENetwork_6_io_to_pes_5_in_valid; // @[pearray.scala 134:13]
  wire [7:0] PENetwork_6_io_to_pes_5_in_bits; // @[pearray.scala 134:13]
  wire  PENetwork_6_io_to_pes_5_out_valid; // @[pearray.scala 134:13]
  wire [7:0] PENetwork_6_io_to_pes_5_out_bits; // @[pearray.scala 134:13]
  wire  PENetwork_6_io_to_pes_6_in_valid; // @[pearray.scala 134:13]
  wire [7:0] PENetwork_6_io_to_pes_6_in_bits; // @[pearray.scala 134:13]
  wire  PENetwork_6_io_to_pes_6_out_valid; // @[pearray.scala 134:13]
  wire [7:0] PENetwork_6_io_to_pes_6_out_bits; // @[pearray.scala 134:13]
  wire  PENetwork_6_io_to_pes_7_in_valid; // @[pearray.scala 134:13]
  wire [7:0] PENetwork_6_io_to_pes_7_in_bits; // @[pearray.scala 134:13]
  wire  PENetwork_6_io_to_pes_7_out_valid; // @[pearray.scala 134:13]
  wire [7:0] PENetwork_6_io_to_pes_7_out_bits; // @[pearray.scala 134:13]
  wire  PENetwork_6_io_to_mem_valid; // @[pearray.scala 134:13]
  wire [7:0] PENetwork_6_io_to_mem_bits; // @[pearray.scala 134:13]
  wire  PENetwork_7_io_to_pes_0_out_valid; // @[pearray.scala 134:13]
  wire [7:0] PENetwork_7_io_to_pes_0_out_bits; // @[pearray.scala 134:13]
  wire  PENetwork_7_io_to_pes_1_in_valid; // @[pearray.scala 134:13]
  wire [7:0] PENetwork_7_io_to_pes_1_in_bits; // @[pearray.scala 134:13]
  wire  PENetwork_7_io_to_pes_1_out_valid; // @[pearray.scala 134:13]
  wire [7:0] PENetwork_7_io_to_pes_1_out_bits; // @[pearray.scala 134:13]
  wire  PENetwork_7_io_to_pes_2_in_valid; // @[pearray.scala 134:13]
  wire [7:0] PENetwork_7_io_to_pes_2_in_bits; // @[pearray.scala 134:13]
  wire  PENetwork_7_io_to_pes_2_out_valid; // @[pearray.scala 134:13]
  wire [7:0] PENetwork_7_io_to_pes_2_out_bits; // @[pearray.scala 134:13]
  wire  PENetwork_7_io_to_pes_3_in_valid; // @[pearray.scala 134:13]
  wire [7:0] PENetwork_7_io_to_pes_3_in_bits; // @[pearray.scala 134:13]
  wire  PENetwork_7_io_to_pes_3_out_valid; // @[pearray.scala 134:13]
  wire [7:0] PENetwork_7_io_to_pes_3_out_bits; // @[pearray.scala 134:13]
  wire  PENetwork_7_io_to_pes_4_in_valid; // @[pearray.scala 134:13]
  wire [7:0] PENetwork_7_io_to_pes_4_in_bits; // @[pearray.scala 134:13]
  wire  PENetwork_7_io_to_pes_4_out_valid; // @[pearray.scala 134:13]
  wire [7:0] PENetwork_7_io_to_pes_4_out_bits; // @[pearray.scala 134:13]
  wire  PENetwork_7_io_to_pes_5_in_valid; // @[pearray.scala 134:13]
  wire [7:0] PENetwork_7_io_to_pes_5_in_bits; // @[pearray.scala 134:13]
  wire  PENetwork_7_io_to_pes_5_out_valid; // @[pearray.scala 134:13]
  wire [7:0] PENetwork_7_io_to_pes_5_out_bits; // @[pearray.scala 134:13]
  wire  PENetwork_7_io_to_pes_6_in_valid; // @[pearray.scala 134:13]
  wire [7:0] PENetwork_7_io_to_pes_6_in_bits; // @[pearray.scala 134:13]
  wire  PENetwork_7_io_to_pes_6_out_valid; // @[pearray.scala 134:13]
  wire [7:0] PENetwork_7_io_to_pes_6_out_bits; // @[pearray.scala 134:13]
  wire  PENetwork_7_io_to_pes_7_in_valid; // @[pearray.scala 134:13]
  wire [7:0] PENetwork_7_io_to_pes_7_in_bits; // @[pearray.scala 134:13]
  wire  PENetwork_7_io_to_pes_7_out_valid; // @[pearray.scala 134:13]
  wire [7:0] PENetwork_7_io_to_pes_7_out_bits; // @[pearray.scala 134:13]
  wire  PENetwork_7_io_to_mem_valid; // @[pearray.scala 134:13]
  wire [7:0] PENetwork_7_io_to_mem_bits; // @[pearray.scala 134:13]
  wire  PENetwork_8_io_to_pes_0_out_valid; // @[pearray.scala 134:13]
  wire [7:0] PENetwork_8_io_to_pes_0_out_bits; // @[pearray.scala 134:13]
  wire  PENetwork_8_io_to_pes_1_in_valid; // @[pearray.scala 134:13]
  wire [7:0] PENetwork_8_io_to_pes_1_in_bits; // @[pearray.scala 134:13]
  wire  PENetwork_8_io_to_pes_1_out_valid; // @[pearray.scala 134:13]
  wire [7:0] PENetwork_8_io_to_pes_1_out_bits; // @[pearray.scala 134:13]
  wire  PENetwork_8_io_to_pes_2_in_valid; // @[pearray.scala 134:13]
  wire [7:0] PENetwork_8_io_to_pes_2_in_bits; // @[pearray.scala 134:13]
  wire  PENetwork_8_io_to_pes_2_out_valid; // @[pearray.scala 134:13]
  wire [7:0] PENetwork_8_io_to_pes_2_out_bits; // @[pearray.scala 134:13]
  wire  PENetwork_8_io_to_pes_3_in_valid; // @[pearray.scala 134:13]
  wire [7:0] PENetwork_8_io_to_pes_3_in_bits; // @[pearray.scala 134:13]
  wire  PENetwork_8_io_to_pes_3_out_valid; // @[pearray.scala 134:13]
  wire [7:0] PENetwork_8_io_to_pes_3_out_bits; // @[pearray.scala 134:13]
  wire  PENetwork_8_io_to_pes_4_in_valid; // @[pearray.scala 134:13]
  wire [7:0] PENetwork_8_io_to_pes_4_in_bits; // @[pearray.scala 134:13]
  wire  PENetwork_8_io_to_pes_4_out_valid; // @[pearray.scala 134:13]
  wire [7:0] PENetwork_8_io_to_pes_4_out_bits; // @[pearray.scala 134:13]
  wire  PENetwork_8_io_to_pes_5_in_valid; // @[pearray.scala 134:13]
  wire [7:0] PENetwork_8_io_to_pes_5_in_bits; // @[pearray.scala 134:13]
  wire  PENetwork_8_io_to_pes_5_out_valid; // @[pearray.scala 134:13]
  wire [7:0] PENetwork_8_io_to_pes_5_out_bits; // @[pearray.scala 134:13]
  wire  PENetwork_8_io_to_pes_6_in_valid; // @[pearray.scala 134:13]
  wire [7:0] PENetwork_8_io_to_pes_6_in_bits; // @[pearray.scala 134:13]
  wire  PENetwork_8_io_to_pes_6_out_valid; // @[pearray.scala 134:13]
  wire [7:0] PENetwork_8_io_to_pes_6_out_bits; // @[pearray.scala 134:13]
  wire  PENetwork_8_io_to_pes_7_in_valid; // @[pearray.scala 134:13]
  wire [7:0] PENetwork_8_io_to_pes_7_in_bits; // @[pearray.scala 134:13]
  wire  PENetwork_8_io_to_pes_7_out_valid; // @[pearray.scala 134:13]
  wire [7:0] PENetwork_8_io_to_pes_7_out_bits; // @[pearray.scala 134:13]
  wire  PENetwork_8_io_to_mem_valid; // @[pearray.scala 134:13]
  wire [7:0] PENetwork_8_io_to_mem_bits; // @[pearray.scala 134:13]
  wire  PENetwork_9_io_to_pes_0_out_valid; // @[pearray.scala 134:13]
  wire [7:0] PENetwork_9_io_to_pes_0_out_bits; // @[pearray.scala 134:13]
  wire  PENetwork_9_io_to_pes_1_in_valid; // @[pearray.scala 134:13]
  wire [7:0] PENetwork_9_io_to_pes_1_in_bits; // @[pearray.scala 134:13]
  wire  PENetwork_9_io_to_pes_1_out_valid; // @[pearray.scala 134:13]
  wire [7:0] PENetwork_9_io_to_pes_1_out_bits; // @[pearray.scala 134:13]
  wire  PENetwork_9_io_to_pes_2_in_valid; // @[pearray.scala 134:13]
  wire [7:0] PENetwork_9_io_to_pes_2_in_bits; // @[pearray.scala 134:13]
  wire  PENetwork_9_io_to_pes_2_out_valid; // @[pearray.scala 134:13]
  wire [7:0] PENetwork_9_io_to_pes_2_out_bits; // @[pearray.scala 134:13]
  wire  PENetwork_9_io_to_pes_3_in_valid; // @[pearray.scala 134:13]
  wire [7:0] PENetwork_9_io_to_pes_3_in_bits; // @[pearray.scala 134:13]
  wire  PENetwork_9_io_to_pes_3_out_valid; // @[pearray.scala 134:13]
  wire [7:0] PENetwork_9_io_to_pes_3_out_bits; // @[pearray.scala 134:13]
  wire  PENetwork_9_io_to_pes_4_in_valid; // @[pearray.scala 134:13]
  wire [7:0] PENetwork_9_io_to_pes_4_in_bits; // @[pearray.scala 134:13]
  wire  PENetwork_9_io_to_pes_4_out_valid; // @[pearray.scala 134:13]
  wire [7:0] PENetwork_9_io_to_pes_4_out_bits; // @[pearray.scala 134:13]
  wire  PENetwork_9_io_to_pes_5_in_valid; // @[pearray.scala 134:13]
  wire [7:0] PENetwork_9_io_to_pes_5_in_bits; // @[pearray.scala 134:13]
  wire  PENetwork_9_io_to_pes_5_out_valid; // @[pearray.scala 134:13]
  wire [7:0] PENetwork_9_io_to_pes_5_out_bits; // @[pearray.scala 134:13]
  wire  PENetwork_9_io_to_pes_6_in_valid; // @[pearray.scala 134:13]
  wire [7:0] PENetwork_9_io_to_pes_6_in_bits; // @[pearray.scala 134:13]
  wire  PENetwork_9_io_to_pes_6_out_valid; // @[pearray.scala 134:13]
  wire [7:0] PENetwork_9_io_to_pes_6_out_bits; // @[pearray.scala 134:13]
  wire  PENetwork_9_io_to_pes_7_in_valid; // @[pearray.scala 134:13]
  wire [7:0] PENetwork_9_io_to_pes_7_in_bits; // @[pearray.scala 134:13]
  wire  PENetwork_9_io_to_pes_7_out_valid; // @[pearray.scala 134:13]
  wire [7:0] PENetwork_9_io_to_pes_7_out_bits; // @[pearray.scala 134:13]
  wire  PENetwork_9_io_to_mem_valid; // @[pearray.scala 134:13]
  wire [7:0] PENetwork_9_io_to_mem_bits; // @[pearray.scala 134:13]
  wire  PENetwork_10_io_to_pes_0_out_valid; // @[pearray.scala 134:13]
  wire [7:0] PENetwork_10_io_to_pes_0_out_bits; // @[pearray.scala 134:13]
  wire  PENetwork_10_io_to_pes_1_in_valid; // @[pearray.scala 134:13]
  wire [7:0] PENetwork_10_io_to_pes_1_in_bits; // @[pearray.scala 134:13]
  wire  PENetwork_10_io_to_pes_1_out_valid; // @[pearray.scala 134:13]
  wire [7:0] PENetwork_10_io_to_pes_1_out_bits; // @[pearray.scala 134:13]
  wire  PENetwork_10_io_to_pes_2_in_valid; // @[pearray.scala 134:13]
  wire [7:0] PENetwork_10_io_to_pes_2_in_bits; // @[pearray.scala 134:13]
  wire  PENetwork_10_io_to_pes_2_out_valid; // @[pearray.scala 134:13]
  wire [7:0] PENetwork_10_io_to_pes_2_out_bits; // @[pearray.scala 134:13]
  wire  PENetwork_10_io_to_pes_3_in_valid; // @[pearray.scala 134:13]
  wire [7:0] PENetwork_10_io_to_pes_3_in_bits; // @[pearray.scala 134:13]
  wire  PENetwork_10_io_to_pes_3_out_valid; // @[pearray.scala 134:13]
  wire [7:0] PENetwork_10_io_to_pes_3_out_bits; // @[pearray.scala 134:13]
  wire  PENetwork_10_io_to_pes_4_in_valid; // @[pearray.scala 134:13]
  wire [7:0] PENetwork_10_io_to_pes_4_in_bits; // @[pearray.scala 134:13]
  wire  PENetwork_10_io_to_pes_4_out_valid; // @[pearray.scala 134:13]
  wire [7:0] PENetwork_10_io_to_pes_4_out_bits; // @[pearray.scala 134:13]
  wire  PENetwork_10_io_to_pes_5_in_valid; // @[pearray.scala 134:13]
  wire [7:0] PENetwork_10_io_to_pes_5_in_bits; // @[pearray.scala 134:13]
  wire  PENetwork_10_io_to_pes_5_out_valid; // @[pearray.scala 134:13]
  wire [7:0] PENetwork_10_io_to_pes_5_out_bits; // @[pearray.scala 134:13]
  wire  PENetwork_10_io_to_pes_6_in_valid; // @[pearray.scala 134:13]
  wire [7:0] PENetwork_10_io_to_pes_6_in_bits; // @[pearray.scala 134:13]
  wire  PENetwork_10_io_to_pes_6_out_valid; // @[pearray.scala 134:13]
  wire [7:0] PENetwork_10_io_to_pes_6_out_bits; // @[pearray.scala 134:13]
  wire  PENetwork_10_io_to_pes_7_in_valid; // @[pearray.scala 134:13]
  wire [7:0] PENetwork_10_io_to_pes_7_in_bits; // @[pearray.scala 134:13]
  wire  PENetwork_10_io_to_pes_7_out_valid; // @[pearray.scala 134:13]
  wire [7:0] PENetwork_10_io_to_pes_7_out_bits; // @[pearray.scala 134:13]
  wire  PENetwork_10_io_to_mem_valid; // @[pearray.scala 134:13]
  wire [7:0] PENetwork_10_io_to_mem_bits; // @[pearray.scala 134:13]
  wire  PENetwork_11_io_to_pes_0_out_valid; // @[pearray.scala 134:13]
  wire [7:0] PENetwork_11_io_to_pes_0_out_bits; // @[pearray.scala 134:13]
  wire  PENetwork_11_io_to_pes_1_in_valid; // @[pearray.scala 134:13]
  wire [7:0] PENetwork_11_io_to_pes_1_in_bits; // @[pearray.scala 134:13]
  wire  PENetwork_11_io_to_pes_1_out_valid; // @[pearray.scala 134:13]
  wire [7:0] PENetwork_11_io_to_pes_1_out_bits; // @[pearray.scala 134:13]
  wire  PENetwork_11_io_to_pes_2_in_valid; // @[pearray.scala 134:13]
  wire [7:0] PENetwork_11_io_to_pes_2_in_bits; // @[pearray.scala 134:13]
  wire  PENetwork_11_io_to_pes_2_out_valid; // @[pearray.scala 134:13]
  wire [7:0] PENetwork_11_io_to_pes_2_out_bits; // @[pearray.scala 134:13]
  wire  PENetwork_11_io_to_pes_3_in_valid; // @[pearray.scala 134:13]
  wire [7:0] PENetwork_11_io_to_pes_3_in_bits; // @[pearray.scala 134:13]
  wire  PENetwork_11_io_to_pes_3_out_valid; // @[pearray.scala 134:13]
  wire [7:0] PENetwork_11_io_to_pes_3_out_bits; // @[pearray.scala 134:13]
  wire  PENetwork_11_io_to_pes_4_in_valid; // @[pearray.scala 134:13]
  wire [7:0] PENetwork_11_io_to_pes_4_in_bits; // @[pearray.scala 134:13]
  wire  PENetwork_11_io_to_pes_4_out_valid; // @[pearray.scala 134:13]
  wire [7:0] PENetwork_11_io_to_pes_4_out_bits; // @[pearray.scala 134:13]
  wire  PENetwork_11_io_to_pes_5_in_valid; // @[pearray.scala 134:13]
  wire [7:0] PENetwork_11_io_to_pes_5_in_bits; // @[pearray.scala 134:13]
  wire  PENetwork_11_io_to_pes_5_out_valid; // @[pearray.scala 134:13]
  wire [7:0] PENetwork_11_io_to_pes_5_out_bits; // @[pearray.scala 134:13]
  wire  PENetwork_11_io_to_pes_6_in_valid; // @[pearray.scala 134:13]
  wire [7:0] PENetwork_11_io_to_pes_6_in_bits; // @[pearray.scala 134:13]
  wire  PENetwork_11_io_to_pes_6_out_valid; // @[pearray.scala 134:13]
  wire [7:0] PENetwork_11_io_to_pes_6_out_bits; // @[pearray.scala 134:13]
  wire  PENetwork_11_io_to_pes_7_in_valid; // @[pearray.scala 134:13]
  wire [7:0] PENetwork_11_io_to_pes_7_in_bits; // @[pearray.scala 134:13]
  wire  PENetwork_11_io_to_pes_7_out_valid; // @[pearray.scala 134:13]
  wire [7:0] PENetwork_11_io_to_pes_7_out_bits; // @[pearray.scala 134:13]
  wire  PENetwork_11_io_to_mem_valid; // @[pearray.scala 134:13]
  wire [7:0] PENetwork_11_io_to_mem_bits; // @[pearray.scala 134:13]
  wire  PENetwork_12_io_to_pes_0_out_valid; // @[pearray.scala 134:13]
  wire [7:0] PENetwork_12_io_to_pes_0_out_bits; // @[pearray.scala 134:13]
  wire  PENetwork_12_io_to_pes_1_in_valid; // @[pearray.scala 134:13]
  wire [7:0] PENetwork_12_io_to_pes_1_in_bits; // @[pearray.scala 134:13]
  wire  PENetwork_12_io_to_pes_1_out_valid; // @[pearray.scala 134:13]
  wire [7:0] PENetwork_12_io_to_pes_1_out_bits; // @[pearray.scala 134:13]
  wire  PENetwork_12_io_to_pes_2_in_valid; // @[pearray.scala 134:13]
  wire [7:0] PENetwork_12_io_to_pes_2_in_bits; // @[pearray.scala 134:13]
  wire  PENetwork_12_io_to_pes_2_out_valid; // @[pearray.scala 134:13]
  wire [7:0] PENetwork_12_io_to_pes_2_out_bits; // @[pearray.scala 134:13]
  wire  PENetwork_12_io_to_pes_3_in_valid; // @[pearray.scala 134:13]
  wire [7:0] PENetwork_12_io_to_pes_3_in_bits; // @[pearray.scala 134:13]
  wire  PENetwork_12_io_to_pes_3_out_valid; // @[pearray.scala 134:13]
  wire [7:0] PENetwork_12_io_to_pes_3_out_bits; // @[pearray.scala 134:13]
  wire  PENetwork_12_io_to_pes_4_in_valid; // @[pearray.scala 134:13]
  wire [7:0] PENetwork_12_io_to_pes_4_in_bits; // @[pearray.scala 134:13]
  wire  PENetwork_12_io_to_pes_4_out_valid; // @[pearray.scala 134:13]
  wire [7:0] PENetwork_12_io_to_pes_4_out_bits; // @[pearray.scala 134:13]
  wire  PENetwork_12_io_to_pes_5_in_valid; // @[pearray.scala 134:13]
  wire [7:0] PENetwork_12_io_to_pes_5_in_bits; // @[pearray.scala 134:13]
  wire  PENetwork_12_io_to_pes_5_out_valid; // @[pearray.scala 134:13]
  wire [7:0] PENetwork_12_io_to_pes_5_out_bits; // @[pearray.scala 134:13]
  wire  PENetwork_12_io_to_pes_6_in_valid; // @[pearray.scala 134:13]
  wire [7:0] PENetwork_12_io_to_pes_6_in_bits; // @[pearray.scala 134:13]
  wire  PENetwork_12_io_to_pes_6_out_valid; // @[pearray.scala 134:13]
  wire [7:0] PENetwork_12_io_to_pes_6_out_bits; // @[pearray.scala 134:13]
  wire  PENetwork_12_io_to_pes_7_in_valid; // @[pearray.scala 134:13]
  wire [7:0] PENetwork_12_io_to_pes_7_in_bits; // @[pearray.scala 134:13]
  wire  PENetwork_12_io_to_pes_7_out_valid; // @[pearray.scala 134:13]
  wire [7:0] PENetwork_12_io_to_pes_7_out_bits; // @[pearray.scala 134:13]
  wire  PENetwork_12_io_to_mem_valid; // @[pearray.scala 134:13]
  wire [7:0] PENetwork_12_io_to_mem_bits; // @[pearray.scala 134:13]
  wire  PENetwork_13_io_to_pes_0_out_valid; // @[pearray.scala 134:13]
  wire [7:0] PENetwork_13_io_to_pes_0_out_bits; // @[pearray.scala 134:13]
  wire  PENetwork_13_io_to_pes_1_in_valid; // @[pearray.scala 134:13]
  wire [7:0] PENetwork_13_io_to_pes_1_in_bits; // @[pearray.scala 134:13]
  wire  PENetwork_13_io_to_pes_1_out_valid; // @[pearray.scala 134:13]
  wire [7:0] PENetwork_13_io_to_pes_1_out_bits; // @[pearray.scala 134:13]
  wire  PENetwork_13_io_to_pes_2_in_valid; // @[pearray.scala 134:13]
  wire [7:0] PENetwork_13_io_to_pes_2_in_bits; // @[pearray.scala 134:13]
  wire  PENetwork_13_io_to_pes_2_out_valid; // @[pearray.scala 134:13]
  wire [7:0] PENetwork_13_io_to_pes_2_out_bits; // @[pearray.scala 134:13]
  wire  PENetwork_13_io_to_pes_3_in_valid; // @[pearray.scala 134:13]
  wire [7:0] PENetwork_13_io_to_pes_3_in_bits; // @[pearray.scala 134:13]
  wire  PENetwork_13_io_to_pes_3_out_valid; // @[pearray.scala 134:13]
  wire [7:0] PENetwork_13_io_to_pes_3_out_bits; // @[pearray.scala 134:13]
  wire  PENetwork_13_io_to_pes_4_in_valid; // @[pearray.scala 134:13]
  wire [7:0] PENetwork_13_io_to_pes_4_in_bits; // @[pearray.scala 134:13]
  wire  PENetwork_13_io_to_pes_4_out_valid; // @[pearray.scala 134:13]
  wire [7:0] PENetwork_13_io_to_pes_4_out_bits; // @[pearray.scala 134:13]
  wire  PENetwork_13_io_to_pes_5_in_valid; // @[pearray.scala 134:13]
  wire [7:0] PENetwork_13_io_to_pes_5_in_bits; // @[pearray.scala 134:13]
  wire  PENetwork_13_io_to_pes_5_out_valid; // @[pearray.scala 134:13]
  wire [7:0] PENetwork_13_io_to_pes_5_out_bits; // @[pearray.scala 134:13]
  wire  PENetwork_13_io_to_pes_6_in_valid; // @[pearray.scala 134:13]
  wire [7:0] PENetwork_13_io_to_pes_6_in_bits; // @[pearray.scala 134:13]
  wire  PENetwork_13_io_to_pes_6_out_valid; // @[pearray.scala 134:13]
  wire [7:0] PENetwork_13_io_to_pes_6_out_bits; // @[pearray.scala 134:13]
  wire  PENetwork_13_io_to_pes_7_in_valid; // @[pearray.scala 134:13]
  wire [7:0] PENetwork_13_io_to_pes_7_in_bits; // @[pearray.scala 134:13]
  wire  PENetwork_13_io_to_pes_7_out_valid; // @[pearray.scala 134:13]
  wire [7:0] PENetwork_13_io_to_pes_7_out_bits; // @[pearray.scala 134:13]
  wire  PENetwork_13_io_to_mem_valid; // @[pearray.scala 134:13]
  wire [7:0] PENetwork_13_io_to_mem_bits; // @[pearray.scala 134:13]
  wire  PENetwork_14_io_to_pes_0_out_valid; // @[pearray.scala 134:13]
  wire [7:0] PENetwork_14_io_to_pes_0_out_bits; // @[pearray.scala 134:13]
  wire  PENetwork_14_io_to_pes_1_in_valid; // @[pearray.scala 134:13]
  wire [7:0] PENetwork_14_io_to_pes_1_in_bits; // @[pearray.scala 134:13]
  wire  PENetwork_14_io_to_pes_1_out_valid; // @[pearray.scala 134:13]
  wire [7:0] PENetwork_14_io_to_pes_1_out_bits; // @[pearray.scala 134:13]
  wire  PENetwork_14_io_to_pes_2_in_valid; // @[pearray.scala 134:13]
  wire [7:0] PENetwork_14_io_to_pes_2_in_bits; // @[pearray.scala 134:13]
  wire  PENetwork_14_io_to_pes_2_out_valid; // @[pearray.scala 134:13]
  wire [7:0] PENetwork_14_io_to_pes_2_out_bits; // @[pearray.scala 134:13]
  wire  PENetwork_14_io_to_pes_3_in_valid; // @[pearray.scala 134:13]
  wire [7:0] PENetwork_14_io_to_pes_3_in_bits; // @[pearray.scala 134:13]
  wire  PENetwork_14_io_to_pes_3_out_valid; // @[pearray.scala 134:13]
  wire [7:0] PENetwork_14_io_to_pes_3_out_bits; // @[pearray.scala 134:13]
  wire  PENetwork_14_io_to_pes_4_in_valid; // @[pearray.scala 134:13]
  wire [7:0] PENetwork_14_io_to_pes_4_in_bits; // @[pearray.scala 134:13]
  wire  PENetwork_14_io_to_pes_4_out_valid; // @[pearray.scala 134:13]
  wire [7:0] PENetwork_14_io_to_pes_4_out_bits; // @[pearray.scala 134:13]
  wire  PENetwork_14_io_to_pes_5_in_valid; // @[pearray.scala 134:13]
  wire [7:0] PENetwork_14_io_to_pes_5_in_bits; // @[pearray.scala 134:13]
  wire  PENetwork_14_io_to_pes_5_out_valid; // @[pearray.scala 134:13]
  wire [7:0] PENetwork_14_io_to_pes_5_out_bits; // @[pearray.scala 134:13]
  wire  PENetwork_14_io_to_pes_6_in_valid; // @[pearray.scala 134:13]
  wire [7:0] PENetwork_14_io_to_pes_6_in_bits; // @[pearray.scala 134:13]
  wire  PENetwork_14_io_to_pes_6_out_valid; // @[pearray.scala 134:13]
  wire [7:0] PENetwork_14_io_to_pes_6_out_bits; // @[pearray.scala 134:13]
  wire  PENetwork_14_io_to_pes_7_in_valid; // @[pearray.scala 134:13]
  wire [7:0] PENetwork_14_io_to_pes_7_in_bits; // @[pearray.scala 134:13]
  wire  PENetwork_14_io_to_pes_7_out_valid; // @[pearray.scala 134:13]
  wire [7:0] PENetwork_14_io_to_pes_7_out_bits; // @[pearray.scala 134:13]
  wire  PENetwork_14_io_to_mem_valid; // @[pearray.scala 134:13]
  wire [7:0] PENetwork_14_io_to_mem_bits; // @[pearray.scala 134:13]
  wire  PENetwork_15_io_to_pes_0_out_valid; // @[pearray.scala 134:13]
  wire [7:0] PENetwork_15_io_to_pes_0_out_bits; // @[pearray.scala 134:13]
  wire  PENetwork_15_io_to_pes_1_in_valid; // @[pearray.scala 134:13]
  wire [7:0] PENetwork_15_io_to_pes_1_in_bits; // @[pearray.scala 134:13]
  wire  PENetwork_15_io_to_pes_1_out_valid; // @[pearray.scala 134:13]
  wire [7:0] PENetwork_15_io_to_pes_1_out_bits; // @[pearray.scala 134:13]
  wire  PENetwork_15_io_to_pes_2_in_valid; // @[pearray.scala 134:13]
  wire [7:0] PENetwork_15_io_to_pes_2_in_bits; // @[pearray.scala 134:13]
  wire  PENetwork_15_io_to_pes_2_out_valid; // @[pearray.scala 134:13]
  wire [7:0] PENetwork_15_io_to_pes_2_out_bits; // @[pearray.scala 134:13]
  wire  PENetwork_15_io_to_pes_3_in_valid; // @[pearray.scala 134:13]
  wire [7:0] PENetwork_15_io_to_pes_3_in_bits; // @[pearray.scala 134:13]
  wire  PENetwork_15_io_to_pes_3_out_valid; // @[pearray.scala 134:13]
  wire [7:0] PENetwork_15_io_to_pes_3_out_bits; // @[pearray.scala 134:13]
  wire  PENetwork_15_io_to_pes_4_in_valid; // @[pearray.scala 134:13]
  wire [7:0] PENetwork_15_io_to_pes_4_in_bits; // @[pearray.scala 134:13]
  wire  PENetwork_15_io_to_pes_4_out_valid; // @[pearray.scala 134:13]
  wire [7:0] PENetwork_15_io_to_pes_4_out_bits; // @[pearray.scala 134:13]
  wire  PENetwork_15_io_to_pes_5_in_valid; // @[pearray.scala 134:13]
  wire [7:0] PENetwork_15_io_to_pes_5_in_bits; // @[pearray.scala 134:13]
  wire  PENetwork_15_io_to_pes_5_out_valid; // @[pearray.scala 134:13]
  wire [7:0] PENetwork_15_io_to_pes_5_out_bits; // @[pearray.scala 134:13]
  wire  PENetwork_15_io_to_pes_6_in_valid; // @[pearray.scala 134:13]
  wire [7:0] PENetwork_15_io_to_pes_6_in_bits; // @[pearray.scala 134:13]
  wire  PENetwork_15_io_to_pes_6_out_valid; // @[pearray.scala 134:13]
  wire [7:0] PENetwork_15_io_to_pes_6_out_bits; // @[pearray.scala 134:13]
  wire  PENetwork_15_io_to_pes_7_in_valid; // @[pearray.scala 134:13]
  wire [7:0] PENetwork_15_io_to_pes_7_in_bits; // @[pearray.scala 134:13]
  wire  PENetwork_15_io_to_pes_7_out_valid; // @[pearray.scala 134:13]
  wire [7:0] PENetwork_15_io_to_pes_7_out_bits; // @[pearray.scala 134:13]
  wire  PENetwork_15_io_to_mem_valid; // @[pearray.scala 134:13]
  wire [7:0] PENetwork_15_io_to_mem_bits; // @[pearray.scala 134:13]
  wire  PENetwork_16_io_to_pes_0_in_valid; // @[pearray.scala 134:13]
  wire [7:0] PENetwork_16_io_to_pes_0_in_bits; // @[pearray.scala 134:13]
  wire  PENetwork_16_io_to_pes_0_out_valid; // @[pearray.scala 134:13]
  wire [7:0] PENetwork_16_io_to_pes_0_out_bits; // @[pearray.scala 134:13]
  wire  PENetwork_16_io_to_pes_1_in_valid; // @[pearray.scala 134:13]
  wire [7:0] PENetwork_16_io_to_pes_1_in_bits; // @[pearray.scala 134:13]
  wire  PENetwork_16_io_to_pes_1_out_valid; // @[pearray.scala 134:13]
  wire [7:0] PENetwork_16_io_to_pes_1_out_bits; // @[pearray.scala 134:13]
  wire  PENetwork_16_io_to_pes_2_in_valid; // @[pearray.scala 134:13]
  wire [7:0] PENetwork_16_io_to_pes_2_in_bits; // @[pearray.scala 134:13]
  wire  PENetwork_16_io_to_pes_2_out_valid; // @[pearray.scala 134:13]
  wire [7:0] PENetwork_16_io_to_pes_2_out_bits; // @[pearray.scala 134:13]
  wire  PENetwork_16_io_to_pes_3_in_valid; // @[pearray.scala 134:13]
  wire [7:0] PENetwork_16_io_to_pes_3_in_bits; // @[pearray.scala 134:13]
  wire  PENetwork_16_io_to_pes_3_out_valid; // @[pearray.scala 134:13]
  wire [7:0] PENetwork_16_io_to_pes_3_out_bits; // @[pearray.scala 134:13]
  wire  PENetwork_16_io_to_pes_4_in_valid; // @[pearray.scala 134:13]
  wire [7:0] PENetwork_16_io_to_pes_4_in_bits; // @[pearray.scala 134:13]
  wire  PENetwork_16_io_to_pes_4_out_valid; // @[pearray.scala 134:13]
  wire [7:0] PENetwork_16_io_to_pes_4_out_bits; // @[pearray.scala 134:13]
  wire  PENetwork_16_io_to_pes_5_in_valid; // @[pearray.scala 134:13]
  wire [7:0] PENetwork_16_io_to_pes_5_in_bits; // @[pearray.scala 134:13]
  wire  PENetwork_16_io_to_pes_5_out_valid; // @[pearray.scala 134:13]
  wire [7:0] PENetwork_16_io_to_pes_5_out_bits; // @[pearray.scala 134:13]
  wire  PENetwork_16_io_to_pes_6_in_valid; // @[pearray.scala 134:13]
  wire [7:0] PENetwork_16_io_to_pes_6_in_bits; // @[pearray.scala 134:13]
  wire  PENetwork_16_io_to_pes_6_out_valid; // @[pearray.scala 134:13]
  wire [7:0] PENetwork_16_io_to_pes_6_out_bits; // @[pearray.scala 134:13]
  wire  PENetwork_16_io_to_pes_7_in_valid; // @[pearray.scala 134:13]
  wire [7:0] PENetwork_16_io_to_pes_7_in_bits; // @[pearray.scala 134:13]
  wire  PENetwork_16_io_to_mem_valid; // @[pearray.scala 134:13]
  wire [7:0] PENetwork_16_io_to_mem_bits; // @[pearray.scala 134:13]
  wire  PENetwork_17_io_to_pes_0_in_valid; // @[pearray.scala 134:13]
  wire [7:0] PENetwork_17_io_to_pes_0_in_bits; // @[pearray.scala 134:13]
  wire  PENetwork_17_io_to_pes_0_out_valid; // @[pearray.scala 134:13]
  wire [7:0] PENetwork_17_io_to_pes_0_out_bits; // @[pearray.scala 134:13]
  wire  PENetwork_17_io_to_pes_1_in_valid; // @[pearray.scala 134:13]
  wire [7:0] PENetwork_17_io_to_pes_1_in_bits; // @[pearray.scala 134:13]
  wire  PENetwork_17_io_to_pes_1_out_valid; // @[pearray.scala 134:13]
  wire [7:0] PENetwork_17_io_to_pes_1_out_bits; // @[pearray.scala 134:13]
  wire  PENetwork_17_io_to_pes_2_in_valid; // @[pearray.scala 134:13]
  wire [7:0] PENetwork_17_io_to_pes_2_in_bits; // @[pearray.scala 134:13]
  wire  PENetwork_17_io_to_pes_2_out_valid; // @[pearray.scala 134:13]
  wire [7:0] PENetwork_17_io_to_pes_2_out_bits; // @[pearray.scala 134:13]
  wire  PENetwork_17_io_to_pes_3_in_valid; // @[pearray.scala 134:13]
  wire [7:0] PENetwork_17_io_to_pes_3_in_bits; // @[pearray.scala 134:13]
  wire  PENetwork_17_io_to_pes_3_out_valid; // @[pearray.scala 134:13]
  wire [7:0] PENetwork_17_io_to_pes_3_out_bits; // @[pearray.scala 134:13]
  wire  PENetwork_17_io_to_pes_4_in_valid; // @[pearray.scala 134:13]
  wire [7:0] PENetwork_17_io_to_pes_4_in_bits; // @[pearray.scala 134:13]
  wire  PENetwork_17_io_to_pes_4_out_valid; // @[pearray.scala 134:13]
  wire [7:0] PENetwork_17_io_to_pes_4_out_bits; // @[pearray.scala 134:13]
  wire  PENetwork_17_io_to_pes_5_in_valid; // @[pearray.scala 134:13]
  wire [7:0] PENetwork_17_io_to_pes_5_in_bits; // @[pearray.scala 134:13]
  wire  PENetwork_17_io_to_pes_5_out_valid; // @[pearray.scala 134:13]
  wire [7:0] PENetwork_17_io_to_pes_5_out_bits; // @[pearray.scala 134:13]
  wire  PENetwork_17_io_to_pes_6_in_valid; // @[pearray.scala 134:13]
  wire [7:0] PENetwork_17_io_to_pes_6_in_bits; // @[pearray.scala 134:13]
  wire  PENetwork_17_io_to_pes_6_out_valid; // @[pearray.scala 134:13]
  wire [7:0] PENetwork_17_io_to_pes_6_out_bits; // @[pearray.scala 134:13]
  wire  PENetwork_17_io_to_pes_7_in_valid; // @[pearray.scala 134:13]
  wire [7:0] PENetwork_17_io_to_pes_7_in_bits; // @[pearray.scala 134:13]
  wire  PENetwork_17_io_to_mem_valid; // @[pearray.scala 134:13]
  wire [7:0] PENetwork_17_io_to_mem_bits; // @[pearray.scala 134:13]
  wire  PENetwork_18_io_to_pes_0_in_valid; // @[pearray.scala 134:13]
  wire [7:0] PENetwork_18_io_to_pes_0_in_bits; // @[pearray.scala 134:13]
  wire  PENetwork_18_io_to_pes_0_out_valid; // @[pearray.scala 134:13]
  wire [7:0] PENetwork_18_io_to_pes_0_out_bits; // @[pearray.scala 134:13]
  wire  PENetwork_18_io_to_pes_1_in_valid; // @[pearray.scala 134:13]
  wire [7:0] PENetwork_18_io_to_pes_1_in_bits; // @[pearray.scala 134:13]
  wire  PENetwork_18_io_to_pes_1_out_valid; // @[pearray.scala 134:13]
  wire [7:0] PENetwork_18_io_to_pes_1_out_bits; // @[pearray.scala 134:13]
  wire  PENetwork_18_io_to_pes_2_in_valid; // @[pearray.scala 134:13]
  wire [7:0] PENetwork_18_io_to_pes_2_in_bits; // @[pearray.scala 134:13]
  wire  PENetwork_18_io_to_pes_2_out_valid; // @[pearray.scala 134:13]
  wire [7:0] PENetwork_18_io_to_pes_2_out_bits; // @[pearray.scala 134:13]
  wire  PENetwork_18_io_to_pes_3_in_valid; // @[pearray.scala 134:13]
  wire [7:0] PENetwork_18_io_to_pes_3_in_bits; // @[pearray.scala 134:13]
  wire  PENetwork_18_io_to_pes_3_out_valid; // @[pearray.scala 134:13]
  wire [7:0] PENetwork_18_io_to_pes_3_out_bits; // @[pearray.scala 134:13]
  wire  PENetwork_18_io_to_pes_4_in_valid; // @[pearray.scala 134:13]
  wire [7:0] PENetwork_18_io_to_pes_4_in_bits; // @[pearray.scala 134:13]
  wire  PENetwork_18_io_to_pes_4_out_valid; // @[pearray.scala 134:13]
  wire [7:0] PENetwork_18_io_to_pes_4_out_bits; // @[pearray.scala 134:13]
  wire  PENetwork_18_io_to_pes_5_in_valid; // @[pearray.scala 134:13]
  wire [7:0] PENetwork_18_io_to_pes_5_in_bits; // @[pearray.scala 134:13]
  wire  PENetwork_18_io_to_pes_5_out_valid; // @[pearray.scala 134:13]
  wire [7:0] PENetwork_18_io_to_pes_5_out_bits; // @[pearray.scala 134:13]
  wire  PENetwork_18_io_to_pes_6_in_valid; // @[pearray.scala 134:13]
  wire [7:0] PENetwork_18_io_to_pes_6_in_bits; // @[pearray.scala 134:13]
  wire  PENetwork_18_io_to_pes_6_out_valid; // @[pearray.scala 134:13]
  wire [7:0] PENetwork_18_io_to_pes_6_out_bits; // @[pearray.scala 134:13]
  wire  PENetwork_18_io_to_pes_7_in_valid; // @[pearray.scala 134:13]
  wire [7:0] PENetwork_18_io_to_pes_7_in_bits; // @[pearray.scala 134:13]
  wire  PENetwork_18_io_to_mem_valid; // @[pearray.scala 134:13]
  wire [7:0] PENetwork_18_io_to_mem_bits; // @[pearray.scala 134:13]
  wire  PENetwork_19_io_to_pes_0_in_valid; // @[pearray.scala 134:13]
  wire [7:0] PENetwork_19_io_to_pes_0_in_bits; // @[pearray.scala 134:13]
  wire  PENetwork_19_io_to_pes_0_out_valid; // @[pearray.scala 134:13]
  wire [7:0] PENetwork_19_io_to_pes_0_out_bits; // @[pearray.scala 134:13]
  wire  PENetwork_19_io_to_pes_1_in_valid; // @[pearray.scala 134:13]
  wire [7:0] PENetwork_19_io_to_pes_1_in_bits; // @[pearray.scala 134:13]
  wire  PENetwork_19_io_to_pes_1_out_valid; // @[pearray.scala 134:13]
  wire [7:0] PENetwork_19_io_to_pes_1_out_bits; // @[pearray.scala 134:13]
  wire  PENetwork_19_io_to_pes_2_in_valid; // @[pearray.scala 134:13]
  wire [7:0] PENetwork_19_io_to_pes_2_in_bits; // @[pearray.scala 134:13]
  wire  PENetwork_19_io_to_pes_2_out_valid; // @[pearray.scala 134:13]
  wire [7:0] PENetwork_19_io_to_pes_2_out_bits; // @[pearray.scala 134:13]
  wire  PENetwork_19_io_to_pes_3_in_valid; // @[pearray.scala 134:13]
  wire [7:0] PENetwork_19_io_to_pes_3_in_bits; // @[pearray.scala 134:13]
  wire  PENetwork_19_io_to_pes_3_out_valid; // @[pearray.scala 134:13]
  wire [7:0] PENetwork_19_io_to_pes_3_out_bits; // @[pearray.scala 134:13]
  wire  PENetwork_19_io_to_pes_4_in_valid; // @[pearray.scala 134:13]
  wire [7:0] PENetwork_19_io_to_pes_4_in_bits; // @[pearray.scala 134:13]
  wire  PENetwork_19_io_to_pes_4_out_valid; // @[pearray.scala 134:13]
  wire [7:0] PENetwork_19_io_to_pes_4_out_bits; // @[pearray.scala 134:13]
  wire  PENetwork_19_io_to_pes_5_in_valid; // @[pearray.scala 134:13]
  wire [7:0] PENetwork_19_io_to_pes_5_in_bits; // @[pearray.scala 134:13]
  wire  PENetwork_19_io_to_pes_5_out_valid; // @[pearray.scala 134:13]
  wire [7:0] PENetwork_19_io_to_pes_5_out_bits; // @[pearray.scala 134:13]
  wire  PENetwork_19_io_to_pes_6_in_valid; // @[pearray.scala 134:13]
  wire [7:0] PENetwork_19_io_to_pes_6_in_bits; // @[pearray.scala 134:13]
  wire  PENetwork_19_io_to_pes_6_out_valid; // @[pearray.scala 134:13]
  wire [7:0] PENetwork_19_io_to_pes_6_out_bits; // @[pearray.scala 134:13]
  wire  PENetwork_19_io_to_pes_7_in_valid; // @[pearray.scala 134:13]
  wire [7:0] PENetwork_19_io_to_pes_7_in_bits; // @[pearray.scala 134:13]
  wire  PENetwork_19_io_to_mem_valid; // @[pearray.scala 134:13]
  wire [7:0] PENetwork_19_io_to_mem_bits; // @[pearray.scala 134:13]
  wire  PENetwork_20_io_to_pes_0_in_valid; // @[pearray.scala 134:13]
  wire [7:0] PENetwork_20_io_to_pes_0_in_bits; // @[pearray.scala 134:13]
  wire  PENetwork_20_io_to_pes_0_out_valid; // @[pearray.scala 134:13]
  wire [7:0] PENetwork_20_io_to_pes_0_out_bits; // @[pearray.scala 134:13]
  wire  PENetwork_20_io_to_pes_1_in_valid; // @[pearray.scala 134:13]
  wire [7:0] PENetwork_20_io_to_pes_1_in_bits; // @[pearray.scala 134:13]
  wire  PENetwork_20_io_to_pes_1_out_valid; // @[pearray.scala 134:13]
  wire [7:0] PENetwork_20_io_to_pes_1_out_bits; // @[pearray.scala 134:13]
  wire  PENetwork_20_io_to_pes_2_in_valid; // @[pearray.scala 134:13]
  wire [7:0] PENetwork_20_io_to_pes_2_in_bits; // @[pearray.scala 134:13]
  wire  PENetwork_20_io_to_pes_2_out_valid; // @[pearray.scala 134:13]
  wire [7:0] PENetwork_20_io_to_pes_2_out_bits; // @[pearray.scala 134:13]
  wire  PENetwork_20_io_to_pes_3_in_valid; // @[pearray.scala 134:13]
  wire [7:0] PENetwork_20_io_to_pes_3_in_bits; // @[pearray.scala 134:13]
  wire  PENetwork_20_io_to_pes_3_out_valid; // @[pearray.scala 134:13]
  wire [7:0] PENetwork_20_io_to_pes_3_out_bits; // @[pearray.scala 134:13]
  wire  PENetwork_20_io_to_pes_4_in_valid; // @[pearray.scala 134:13]
  wire [7:0] PENetwork_20_io_to_pes_4_in_bits; // @[pearray.scala 134:13]
  wire  PENetwork_20_io_to_pes_4_out_valid; // @[pearray.scala 134:13]
  wire [7:0] PENetwork_20_io_to_pes_4_out_bits; // @[pearray.scala 134:13]
  wire  PENetwork_20_io_to_pes_5_in_valid; // @[pearray.scala 134:13]
  wire [7:0] PENetwork_20_io_to_pes_5_in_bits; // @[pearray.scala 134:13]
  wire  PENetwork_20_io_to_pes_5_out_valid; // @[pearray.scala 134:13]
  wire [7:0] PENetwork_20_io_to_pes_5_out_bits; // @[pearray.scala 134:13]
  wire  PENetwork_20_io_to_pes_6_in_valid; // @[pearray.scala 134:13]
  wire [7:0] PENetwork_20_io_to_pes_6_in_bits; // @[pearray.scala 134:13]
  wire  PENetwork_20_io_to_pes_6_out_valid; // @[pearray.scala 134:13]
  wire [7:0] PENetwork_20_io_to_pes_6_out_bits; // @[pearray.scala 134:13]
  wire  PENetwork_20_io_to_pes_7_in_valid; // @[pearray.scala 134:13]
  wire [7:0] PENetwork_20_io_to_pes_7_in_bits; // @[pearray.scala 134:13]
  wire  PENetwork_20_io_to_mem_valid; // @[pearray.scala 134:13]
  wire [7:0] PENetwork_20_io_to_mem_bits; // @[pearray.scala 134:13]
  wire  PENetwork_21_io_to_pes_0_in_valid; // @[pearray.scala 134:13]
  wire [7:0] PENetwork_21_io_to_pes_0_in_bits; // @[pearray.scala 134:13]
  wire  PENetwork_21_io_to_pes_0_out_valid; // @[pearray.scala 134:13]
  wire [7:0] PENetwork_21_io_to_pes_0_out_bits; // @[pearray.scala 134:13]
  wire  PENetwork_21_io_to_pes_1_in_valid; // @[pearray.scala 134:13]
  wire [7:0] PENetwork_21_io_to_pes_1_in_bits; // @[pearray.scala 134:13]
  wire  PENetwork_21_io_to_pes_1_out_valid; // @[pearray.scala 134:13]
  wire [7:0] PENetwork_21_io_to_pes_1_out_bits; // @[pearray.scala 134:13]
  wire  PENetwork_21_io_to_pes_2_in_valid; // @[pearray.scala 134:13]
  wire [7:0] PENetwork_21_io_to_pes_2_in_bits; // @[pearray.scala 134:13]
  wire  PENetwork_21_io_to_pes_2_out_valid; // @[pearray.scala 134:13]
  wire [7:0] PENetwork_21_io_to_pes_2_out_bits; // @[pearray.scala 134:13]
  wire  PENetwork_21_io_to_pes_3_in_valid; // @[pearray.scala 134:13]
  wire [7:0] PENetwork_21_io_to_pes_3_in_bits; // @[pearray.scala 134:13]
  wire  PENetwork_21_io_to_pes_3_out_valid; // @[pearray.scala 134:13]
  wire [7:0] PENetwork_21_io_to_pes_3_out_bits; // @[pearray.scala 134:13]
  wire  PENetwork_21_io_to_pes_4_in_valid; // @[pearray.scala 134:13]
  wire [7:0] PENetwork_21_io_to_pes_4_in_bits; // @[pearray.scala 134:13]
  wire  PENetwork_21_io_to_pes_4_out_valid; // @[pearray.scala 134:13]
  wire [7:0] PENetwork_21_io_to_pes_4_out_bits; // @[pearray.scala 134:13]
  wire  PENetwork_21_io_to_pes_5_in_valid; // @[pearray.scala 134:13]
  wire [7:0] PENetwork_21_io_to_pes_5_in_bits; // @[pearray.scala 134:13]
  wire  PENetwork_21_io_to_pes_5_out_valid; // @[pearray.scala 134:13]
  wire [7:0] PENetwork_21_io_to_pes_5_out_bits; // @[pearray.scala 134:13]
  wire  PENetwork_21_io_to_pes_6_in_valid; // @[pearray.scala 134:13]
  wire [7:0] PENetwork_21_io_to_pes_6_in_bits; // @[pearray.scala 134:13]
  wire  PENetwork_21_io_to_pes_6_out_valid; // @[pearray.scala 134:13]
  wire [7:0] PENetwork_21_io_to_pes_6_out_bits; // @[pearray.scala 134:13]
  wire  PENetwork_21_io_to_pes_7_in_valid; // @[pearray.scala 134:13]
  wire [7:0] PENetwork_21_io_to_pes_7_in_bits; // @[pearray.scala 134:13]
  wire  PENetwork_21_io_to_mem_valid; // @[pearray.scala 134:13]
  wire [7:0] PENetwork_21_io_to_mem_bits; // @[pearray.scala 134:13]
  wire  PENetwork_22_io_to_pes_0_in_valid; // @[pearray.scala 134:13]
  wire [7:0] PENetwork_22_io_to_pes_0_in_bits; // @[pearray.scala 134:13]
  wire  PENetwork_22_io_to_pes_0_out_valid; // @[pearray.scala 134:13]
  wire [7:0] PENetwork_22_io_to_pes_0_out_bits; // @[pearray.scala 134:13]
  wire  PENetwork_22_io_to_pes_1_in_valid; // @[pearray.scala 134:13]
  wire [7:0] PENetwork_22_io_to_pes_1_in_bits; // @[pearray.scala 134:13]
  wire  PENetwork_22_io_to_pes_1_out_valid; // @[pearray.scala 134:13]
  wire [7:0] PENetwork_22_io_to_pes_1_out_bits; // @[pearray.scala 134:13]
  wire  PENetwork_22_io_to_pes_2_in_valid; // @[pearray.scala 134:13]
  wire [7:0] PENetwork_22_io_to_pes_2_in_bits; // @[pearray.scala 134:13]
  wire  PENetwork_22_io_to_pes_2_out_valid; // @[pearray.scala 134:13]
  wire [7:0] PENetwork_22_io_to_pes_2_out_bits; // @[pearray.scala 134:13]
  wire  PENetwork_22_io_to_pes_3_in_valid; // @[pearray.scala 134:13]
  wire [7:0] PENetwork_22_io_to_pes_3_in_bits; // @[pearray.scala 134:13]
  wire  PENetwork_22_io_to_pes_3_out_valid; // @[pearray.scala 134:13]
  wire [7:0] PENetwork_22_io_to_pes_3_out_bits; // @[pearray.scala 134:13]
  wire  PENetwork_22_io_to_pes_4_in_valid; // @[pearray.scala 134:13]
  wire [7:0] PENetwork_22_io_to_pes_4_in_bits; // @[pearray.scala 134:13]
  wire  PENetwork_22_io_to_pes_4_out_valid; // @[pearray.scala 134:13]
  wire [7:0] PENetwork_22_io_to_pes_4_out_bits; // @[pearray.scala 134:13]
  wire  PENetwork_22_io_to_pes_5_in_valid; // @[pearray.scala 134:13]
  wire [7:0] PENetwork_22_io_to_pes_5_in_bits; // @[pearray.scala 134:13]
  wire  PENetwork_22_io_to_pes_5_out_valid; // @[pearray.scala 134:13]
  wire [7:0] PENetwork_22_io_to_pes_5_out_bits; // @[pearray.scala 134:13]
  wire  PENetwork_22_io_to_pes_6_in_valid; // @[pearray.scala 134:13]
  wire [7:0] PENetwork_22_io_to_pes_6_in_bits; // @[pearray.scala 134:13]
  wire  PENetwork_22_io_to_pes_6_out_valid; // @[pearray.scala 134:13]
  wire [7:0] PENetwork_22_io_to_pes_6_out_bits; // @[pearray.scala 134:13]
  wire  PENetwork_22_io_to_pes_7_in_valid; // @[pearray.scala 134:13]
  wire [7:0] PENetwork_22_io_to_pes_7_in_bits; // @[pearray.scala 134:13]
  wire  PENetwork_22_io_to_mem_valid; // @[pearray.scala 134:13]
  wire [7:0] PENetwork_22_io_to_mem_bits; // @[pearray.scala 134:13]
  wire  PENetwork_23_io_to_pes_0_in_valid; // @[pearray.scala 134:13]
  wire [7:0] PENetwork_23_io_to_pes_0_in_bits; // @[pearray.scala 134:13]
  wire  PENetwork_23_io_to_pes_0_out_valid; // @[pearray.scala 134:13]
  wire [7:0] PENetwork_23_io_to_pes_0_out_bits; // @[pearray.scala 134:13]
  wire  PENetwork_23_io_to_pes_1_in_valid; // @[pearray.scala 134:13]
  wire [7:0] PENetwork_23_io_to_pes_1_in_bits; // @[pearray.scala 134:13]
  wire  PENetwork_23_io_to_pes_1_out_valid; // @[pearray.scala 134:13]
  wire [7:0] PENetwork_23_io_to_pes_1_out_bits; // @[pearray.scala 134:13]
  wire  PENetwork_23_io_to_pes_2_in_valid; // @[pearray.scala 134:13]
  wire [7:0] PENetwork_23_io_to_pes_2_in_bits; // @[pearray.scala 134:13]
  wire  PENetwork_23_io_to_pes_2_out_valid; // @[pearray.scala 134:13]
  wire [7:0] PENetwork_23_io_to_pes_2_out_bits; // @[pearray.scala 134:13]
  wire  PENetwork_23_io_to_pes_3_in_valid; // @[pearray.scala 134:13]
  wire [7:0] PENetwork_23_io_to_pes_3_in_bits; // @[pearray.scala 134:13]
  wire  PENetwork_23_io_to_pes_3_out_valid; // @[pearray.scala 134:13]
  wire [7:0] PENetwork_23_io_to_pes_3_out_bits; // @[pearray.scala 134:13]
  wire  PENetwork_23_io_to_pes_4_in_valid; // @[pearray.scala 134:13]
  wire [7:0] PENetwork_23_io_to_pes_4_in_bits; // @[pearray.scala 134:13]
  wire  PENetwork_23_io_to_pes_4_out_valid; // @[pearray.scala 134:13]
  wire [7:0] PENetwork_23_io_to_pes_4_out_bits; // @[pearray.scala 134:13]
  wire  PENetwork_23_io_to_pes_5_in_valid; // @[pearray.scala 134:13]
  wire [7:0] PENetwork_23_io_to_pes_5_in_bits; // @[pearray.scala 134:13]
  wire  PENetwork_23_io_to_pes_5_out_valid; // @[pearray.scala 134:13]
  wire [7:0] PENetwork_23_io_to_pes_5_out_bits; // @[pearray.scala 134:13]
  wire  PENetwork_23_io_to_pes_6_in_valid; // @[pearray.scala 134:13]
  wire [7:0] PENetwork_23_io_to_pes_6_in_bits; // @[pearray.scala 134:13]
  wire  PENetwork_23_io_to_pes_6_out_valid; // @[pearray.scala 134:13]
  wire [7:0] PENetwork_23_io_to_pes_6_out_bits; // @[pearray.scala 134:13]
  wire  PENetwork_23_io_to_pes_7_in_valid; // @[pearray.scala 134:13]
  wire [7:0] PENetwork_23_io_to_pes_7_in_bits; // @[pearray.scala 134:13]
  wire  PENetwork_23_io_to_mem_valid; // @[pearray.scala 134:13]
  wire [7:0] PENetwork_23_io_to_mem_bits; // @[pearray.scala 134:13]
  wire  PENetwork_24_io_to_pes_0_in_valid; // @[pearray.scala 134:13]
  wire [7:0] PENetwork_24_io_to_pes_0_in_bits; // @[pearray.scala 134:13]
  wire  PENetwork_24_io_to_pes_0_out_valid; // @[pearray.scala 134:13]
  wire [7:0] PENetwork_24_io_to_pes_0_out_bits; // @[pearray.scala 134:13]
  wire  PENetwork_24_io_to_pes_1_in_valid; // @[pearray.scala 134:13]
  wire [7:0] PENetwork_24_io_to_pes_1_in_bits; // @[pearray.scala 134:13]
  wire  PENetwork_24_io_to_pes_1_out_valid; // @[pearray.scala 134:13]
  wire [7:0] PENetwork_24_io_to_pes_1_out_bits; // @[pearray.scala 134:13]
  wire  PENetwork_24_io_to_pes_2_in_valid; // @[pearray.scala 134:13]
  wire [7:0] PENetwork_24_io_to_pes_2_in_bits; // @[pearray.scala 134:13]
  wire  PENetwork_24_io_to_pes_2_out_valid; // @[pearray.scala 134:13]
  wire [7:0] PENetwork_24_io_to_pes_2_out_bits; // @[pearray.scala 134:13]
  wire  PENetwork_24_io_to_pes_3_in_valid; // @[pearray.scala 134:13]
  wire [7:0] PENetwork_24_io_to_pes_3_in_bits; // @[pearray.scala 134:13]
  wire  PENetwork_24_io_to_pes_3_out_valid; // @[pearray.scala 134:13]
  wire [7:0] PENetwork_24_io_to_pes_3_out_bits; // @[pearray.scala 134:13]
  wire  PENetwork_24_io_to_pes_4_in_valid; // @[pearray.scala 134:13]
  wire [7:0] PENetwork_24_io_to_pes_4_in_bits; // @[pearray.scala 134:13]
  wire  PENetwork_24_io_to_pes_4_out_valid; // @[pearray.scala 134:13]
  wire [7:0] PENetwork_24_io_to_pes_4_out_bits; // @[pearray.scala 134:13]
  wire  PENetwork_24_io_to_pes_5_in_valid; // @[pearray.scala 134:13]
  wire [7:0] PENetwork_24_io_to_pes_5_in_bits; // @[pearray.scala 134:13]
  wire  PENetwork_24_io_to_pes_5_out_valid; // @[pearray.scala 134:13]
  wire [7:0] PENetwork_24_io_to_pes_5_out_bits; // @[pearray.scala 134:13]
  wire  PENetwork_24_io_to_pes_6_in_valid; // @[pearray.scala 134:13]
  wire [7:0] PENetwork_24_io_to_pes_6_in_bits; // @[pearray.scala 134:13]
  wire  PENetwork_24_io_to_pes_6_out_valid; // @[pearray.scala 134:13]
  wire [7:0] PENetwork_24_io_to_pes_6_out_bits; // @[pearray.scala 134:13]
  wire  PENetwork_24_io_to_pes_7_in_valid; // @[pearray.scala 134:13]
  wire [7:0] PENetwork_24_io_to_pes_7_in_bits; // @[pearray.scala 134:13]
  wire  PENetwork_24_io_to_mem_valid; // @[pearray.scala 134:13]
  wire [7:0] PENetwork_24_io_to_mem_bits; // @[pearray.scala 134:13]
  wire  PENetwork_25_io_to_pes_0_in_valid; // @[pearray.scala 134:13]
  wire [7:0] PENetwork_25_io_to_pes_0_in_bits; // @[pearray.scala 134:13]
  wire  PENetwork_25_io_to_pes_0_out_valid; // @[pearray.scala 134:13]
  wire [7:0] PENetwork_25_io_to_pes_0_out_bits; // @[pearray.scala 134:13]
  wire  PENetwork_25_io_to_pes_1_in_valid; // @[pearray.scala 134:13]
  wire [7:0] PENetwork_25_io_to_pes_1_in_bits; // @[pearray.scala 134:13]
  wire  PENetwork_25_io_to_pes_1_out_valid; // @[pearray.scala 134:13]
  wire [7:0] PENetwork_25_io_to_pes_1_out_bits; // @[pearray.scala 134:13]
  wire  PENetwork_25_io_to_pes_2_in_valid; // @[pearray.scala 134:13]
  wire [7:0] PENetwork_25_io_to_pes_2_in_bits; // @[pearray.scala 134:13]
  wire  PENetwork_25_io_to_pes_2_out_valid; // @[pearray.scala 134:13]
  wire [7:0] PENetwork_25_io_to_pes_2_out_bits; // @[pearray.scala 134:13]
  wire  PENetwork_25_io_to_pes_3_in_valid; // @[pearray.scala 134:13]
  wire [7:0] PENetwork_25_io_to_pes_3_in_bits; // @[pearray.scala 134:13]
  wire  PENetwork_25_io_to_pes_3_out_valid; // @[pearray.scala 134:13]
  wire [7:0] PENetwork_25_io_to_pes_3_out_bits; // @[pearray.scala 134:13]
  wire  PENetwork_25_io_to_pes_4_in_valid; // @[pearray.scala 134:13]
  wire [7:0] PENetwork_25_io_to_pes_4_in_bits; // @[pearray.scala 134:13]
  wire  PENetwork_25_io_to_pes_4_out_valid; // @[pearray.scala 134:13]
  wire [7:0] PENetwork_25_io_to_pes_4_out_bits; // @[pearray.scala 134:13]
  wire  PENetwork_25_io_to_pes_5_in_valid; // @[pearray.scala 134:13]
  wire [7:0] PENetwork_25_io_to_pes_5_in_bits; // @[pearray.scala 134:13]
  wire  PENetwork_25_io_to_pes_5_out_valid; // @[pearray.scala 134:13]
  wire [7:0] PENetwork_25_io_to_pes_5_out_bits; // @[pearray.scala 134:13]
  wire  PENetwork_25_io_to_pes_6_in_valid; // @[pearray.scala 134:13]
  wire [7:0] PENetwork_25_io_to_pes_6_in_bits; // @[pearray.scala 134:13]
  wire  PENetwork_25_io_to_pes_6_out_valid; // @[pearray.scala 134:13]
  wire [7:0] PENetwork_25_io_to_pes_6_out_bits; // @[pearray.scala 134:13]
  wire  PENetwork_25_io_to_pes_7_in_valid; // @[pearray.scala 134:13]
  wire [7:0] PENetwork_25_io_to_pes_7_in_bits; // @[pearray.scala 134:13]
  wire  PENetwork_25_io_to_mem_valid; // @[pearray.scala 134:13]
  wire [7:0] PENetwork_25_io_to_mem_bits; // @[pearray.scala 134:13]
  wire  PENetwork_26_io_to_pes_0_in_valid; // @[pearray.scala 134:13]
  wire [7:0] PENetwork_26_io_to_pes_0_in_bits; // @[pearray.scala 134:13]
  wire  PENetwork_26_io_to_pes_0_out_valid; // @[pearray.scala 134:13]
  wire [7:0] PENetwork_26_io_to_pes_0_out_bits; // @[pearray.scala 134:13]
  wire  PENetwork_26_io_to_pes_1_in_valid; // @[pearray.scala 134:13]
  wire [7:0] PENetwork_26_io_to_pes_1_in_bits; // @[pearray.scala 134:13]
  wire  PENetwork_26_io_to_pes_1_out_valid; // @[pearray.scala 134:13]
  wire [7:0] PENetwork_26_io_to_pes_1_out_bits; // @[pearray.scala 134:13]
  wire  PENetwork_26_io_to_pes_2_in_valid; // @[pearray.scala 134:13]
  wire [7:0] PENetwork_26_io_to_pes_2_in_bits; // @[pearray.scala 134:13]
  wire  PENetwork_26_io_to_pes_2_out_valid; // @[pearray.scala 134:13]
  wire [7:0] PENetwork_26_io_to_pes_2_out_bits; // @[pearray.scala 134:13]
  wire  PENetwork_26_io_to_pes_3_in_valid; // @[pearray.scala 134:13]
  wire [7:0] PENetwork_26_io_to_pes_3_in_bits; // @[pearray.scala 134:13]
  wire  PENetwork_26_io_to_pes_3_out_valid; // @[pearray.scala 134:13]
  wire [7:0] PENetwork_26_io_to_pes_3_out_bits; // @[pearray.scala 134:13]
  wire  PENetwork_26_io_to_pes_4_in_valid; // @[pearray.scala 134:13]
  wire [7:0] PENetwork_26_io_to_pes_4_in_bits; // @[pearray.scala 134:13]
  wire  PENetwork_26_io_to_pes_4_out_valid; // @[pearray.scala 134:13]
  wire [7:0] PENetwork_26_io_to_pes_4_out_bits; // @[pearray.scala 134:13]
  wire  PENetwork_26_io_to_pes_5_in_valid; // @[pearray.scala 134:13]
  wire [7:0] PENetwork_26_io_to_pes_5_in_bits; // @[pearray.scala 134:13]
  wire  PENetwork_26_io_to_pes_5_out_valid; // @[pearray.scala 134:13]
  wire [7:0] PENetwork_26_io_to_pes_5_out_bits; // @[pearray.scala 134:13]
  wire  PENetwork_26_io_to_pes_6_in_valid; // @[pearray.scala 134:13]
  wire [7:0] PENetwork_26_io_to_pes_6_in_bits; // @[pearray.scala 134:13]
  wire  PENetwork_26_io_to_pes_6_out_valid; // @[pearray.scala 134:13]
  wire [7:0] PENetwork_26_io_to_pes_6_out_bits; // @[pearray.scala 134:13]
  wire  PENetwork_26_io_to_pes_7_in_valid; // @[pearray.scala 134:13]
  wire [7:0] PENetwork_26_io_to_pes_7_in_bits; // @[pearray.scala 134:13]
  wire  PENetwork_26_io_to_mem_valid; // @[pearray.scala 134:13]
  wire [7:0] PENetwork_26_io_to_mem_bits; // @[pearray.scala 134:13]
  wire  PENetwork_27_io_to_pes_0_in_valid; // @[pearray.scala 134:13]
  wire [7:0] PENetwork_27_io_to_pes_0_in_bits; // @[pearray.scala 134:13]
  wire  PENetwork_27_io_to_pes_0_out_valid; // @[pearray.scala 134:13]
  wire [7:0] PENetwork_27_io_to_pes_0_out_bits; // @[pearray.scala 134:13]
  wire  PENetwork_27_io_to_pes_1_in_valid; // @[pearray.scala 134:13]
  wire [7:0] PENetwork_27_io_to_pes_1_in_bits; // @[pearray.scala 134:13]
  wire  PENetwork_27_io_to_pes_1_out_valid; // @[pearray.scala 134:13]
  wire [7:0] PENetwork_27_io_to_pes_1_out_bits; // @[pearray.scala 134:13]
  wire  PENetwork_27_io_to_pes_2_in_valid; // @[pearray.scala 134:13]
  wire [7:0] PENetwork_27_io_to_pes_2_in_bits; // @[pearray.scala 134:13]
  wire  PENetwork_27_io_to_pes_2_out_valid; // @[pearray.scala 134:13]
  wire [7:0] PENetwork_27_io_to_pes_2_out_bits; // @[pearray.scala 134:13]
  wire  PENetwork_27_io_to_pes_3_in_valid; // @[pearray.scala 134:13]
  wire [7:0] PENetwork_27_io_to_pes_3_in_bits; // @[pearray.scala 134:13]
  wire  PENetwork_27_io_to_pes_3_out_valid; // @[pearray.scala 134:13]
  wire [7:0] PENetwork_27_io_to_pes_3_out_bits; // @[pearray.scala 134:13]
  wire  PENetwork_27_io_to_pes_4_in_valid; // @[pearray.scala 134:13]
  wire [7:0] PENetwork_27_io_to_pes_4_in_bits; // @[pearray.scala 134:13]
  wire  PENetwork_27_io_to_pes_4_out_valid; // @[pearray.scala 134:13]
  wire [7:0] PENetwork_27_io_to_pes_4_out_bits; // @[pearray.scala 134:13]
  wire  PENetwork_27_io_to_pes_5_in_valid; // @[pearray.scala 134:13]
  wire [7:0] PENetwork_27_io_to_pes_5_in_bits; // @[pearray.scala 134:13]
  wire  PENetwork_27_io_to_pes_5_out_valid; // @[pearray.scala 134:13]
  wire [7:0] PENetwork_27_io_to_pes_5_out_bits; // @[pearray.scala 134:13]
  wire  PENetwork_27_io_to_pes_6_in_valid; // @[pearray.scala 134:13]
  wire [7:0] PENetwork_27_io_to_pes_6_in_bits; // @[pearray.scala 134:13]
  wire  PENetwork_27_io_to_pes_6_out_valid; // @[pearray.scala 134:13]
  wire [7:0] PENetwork_27_io_to_pes_6_out_bits; // @[pearray.scala 134:13]
  wire  PENetwork_27_io_to_pes_7_in_valid; // @[pearray.scala 134:13]
  wire [7:0] PENetwork_27_io_to_pes_7_in_bits; // @[pearray.scala 134:13]
  wire  PENetwork_27_io_to_mem_valid; // @[pearray.scala 134:13]
  wire [7:0] PENetwork_27_io_to_mem_bits; // @[pearray.scala 134:13]
  wire  PENetwork_28_io_to_pes_0_in_valid; // @[pearray.scala 134:13]
  wire [7:0] PENetwork_28_io_to_pes_0_in_bits; // @[pearray.scala 134:13]
  wire  PENetwork_28_io_to_pes_0_out_valid; // @[pearray.scala 134:13]
  wire [7:0] PENetwork_28_io_to_pes_0_out_bits; // @[pearray.scala 134:13]
  wire  PENetwork_28_io_to_pes_1_in_valid; // @[pearray.scala 134:13]
  wire [7:0] PENetwork_28_io_to_pes_1_in_bits; // @[pearray.scala 134:13]
  wire  PENetwork_28_io_to_pes_1_out_valid; // @[pearray.scala 134:13]
  wire [7:0] PENetwork_28_io_to_pes_1_out_bits; // @[pearray.scala 134:13]
  wire  PENetwork_28_io_to_pes_2_in_valid; // @[pearray.scala 134:13]
  wire [7:0] PENetwork_28_io_to_pes_2_in_bits; // @[pearray.scala 134:13]
  wire  PENetwork_28_io_to_pes_2_out_valid; // @[pearray.scala 134:13]
  wire [7:0] PENetwork_28_io_to_pes_2_out_bits; // @[pearray.scala 134:13]
  wire  PENetwork_28_io_to_pes_3_in_valid; // @[pearray.scala 134:13]
  wire [7:0] PENetwork_28_io_to_pes_3_in_bits; // @[pearray.scala 134:13]
  wire  PENetwork_28_io_to_pes_3_out_valid; // @[pearray.scala 134:13]
  wire [7:0] PENetwork_28_io_to_pes_3_out_bits; // @[pearray.scala 134:13]
  wire  PENetwork_28_io_to_pes_4_in_valid; // @[pearray.scala 134:13]
  wire [7:0] PENetwork_28_io_to_pes_4_in_bits; // @[pearray.scala 134:13]
  wire  PENetwork_28_io_to_pes_4_out_valid; // @[pearray.scala 134:13]
  wire [7:0] PENetwork_28_io_to_pes_4_out_bits; // @[pearray.scala 134:13]
  wire  PENetwork_28_io_to_pes_5_in_valid; // @[pearray.scala 134:13]
  wire [7:0] PENetwork_28_io_to_pes_5_in_bits; // @[pearray.scala 134:13]
  wire  PENetwork_28_io_to_pes_5_out_valid; // @[pearray.scala 134:13]
  wire [7:0] PENetwork_28_io_to_pes_5_out_bits; // @[pearray.scala 134:13]
  wire  PENetwork_28_io_to_pes_6_in_valid; // @[pearray.scala 134:13]
  wire [7:0] PENetwork_28_io_to_pes_6_in_bits; // @[pearray.scala 134:13]
  wire  PENetwork_28_io_to_pes_6_out_valid; // @[pearray.scala 134:13]
  wire [7:0] PENetwork_28_io_to_pes_6_out_bits; // @[pearray.scala 134:13]
  wire  PENetwork_28_io_to_pes_7_in_valid; // @[pearray.scala 134:13]
  wire [7:0] PENetwork_28_io_to_pes_7_in_bits; // @[pearray.scala 134:13]
  wire  PENetwork_28_io_to_mem_valid; // @[pearray.scala 134:13]
  wire [7:0] PENetwork_28_io_to_mem_bits; // @[pearray.scala 134:13]
  wire  PENetwork_29_io_to_pes_0_in_valid; // @[pearray.scala 134:13]
  wire [7:0] PENetwork_29_io_to_pes_0_in_bits; // @[pearray.scala 134:13]
  wire  PENetwork_29_io_to_pes_0_out_valid; // @[pearray.scala 134:13]
  wire [7:0] PENetwork_29_io_to_pes_0_out_bits; // @[pearray.scala 134:13]
  wire  PENetwork_29_io_to_pes_1_in_valid; // @[pearray.scala 134:13]
  wire [7:0] PENetwork_29_io_to_pes_1_in_bits; // @[pearray.scala 134:13]
  wire  PENetwork_29_io_to_pes_1_out_valid; // @[pearray.scala 134:13]
  wire [7:0] PENetwork_29_io_to_pes_1_out_bits; // @[pearray.scala 134:13]
  wire  PENetwork_29_io_to_pes_2_in_valid; // @[pearray.scala 134:13]
  wire [7:0] PENetwork_29_io_to_pes_2_in_bits; // @[pearray.scala 134:13]
  wire  PENetwork_29_io_to_pes_2_out_valid; // @[pearray.scala 134:13]
  wire [7:0] PENetwork_29_io_to_pes_2_out_bits; // @[pearray.scala 134:13]
  wire  PENetwork_29_io_to_pes_3_in_valid; // @[pearray.scala 134:13]
  wire [7:0] PENetwork_29_io_to_pes_3_in_bits; // @[pearray.scala 134:13]
  wire  PENetwork_29_io_to_pes_3_out_valid; // @[pearray.scala 134:13]
  wire [7:0] PENetwork_29_io_to_pes_3_out_bits; // @[pearray.scala 134:13]
  wire  PENetwork_29_io_to_pes_4_in_valid; // @[pearray.scala 134:13]
  wire [7:0] PENetwork_29_io_to_pes_4_in_bits; // @[pearray.scala 134:13]
  wire  PENetwork_29_io_to_pes_4_out_valid; // @[pearray.scala 134:13]
  wire [7:0] PENetwork_29_io_to_pes_4_out_bits; // @[pearray.scala 134:13]
  wire  PENetwork_29_io_to_pes_5_in_valid; // @[pearray.scala 134:13]
  wire [7:0] PENetwork_29_io_to_pes_5_in_bits; // @[pearray.scala 134:13]
  wire  PENetwork_29_io_to_pes_5_out_valid; // @[pearray.scala 134:13]
  wire [7:0] PENetwork_29_io_to_pes_5_out_bits; // @[pearray.scala 134:13]
  wire  PENetwork_29_io_to_pes_6_in_valid; // @[pearray.scala 134:13]
  wire [7:0] PENetwork_29_io_to_pes_6_in_bits; // @[pearray.scala 134:13]
  wire  PENetwork_29_io_to_pes_6_out_valid; // @[pearray.scala 134:13]
  wire [7:0] PENetwork_29_io_to_pes_6_out_bits; // @[pearray.scala 134:13]
  wire  PENetwork_29_io_to_pes_7_in_valid; // @[pearray.scala 134:13]
  wire [7:0] PENetwork_29_io_to_pes_7_in_bits; // @[pearray.scala 134:13]
  wire  PENetwork_29_io_to_mem_valid; // @[pearray.scala 134:13]
  wire [7:0] PENetwork_29_io_to_mem_bits; // @[pearray.scala 134:13]
  wire  PENetwork_30_io_to_pes_0_in_valid; // @[pearray.scala 134:13]
  wire [7:0] PENetwork_30_io_to_pes_0_in_bits; // @[pearray.scala 134:13]
  wire  PENetwork_30_io_to_pes_0_out_valid; // @[pearray.scala 134:13]
  wire [7:0] PENetwork_30_io_to_pes_0_out_bits; // @[pearray.scala 134:13]
  wire  PENetwork_30_io_to_pes_1_in_valid; // @[pearray.scala 134:13]
  wire [7:0] PENetwork_30_io_to_pes_1_in_bits; // @[pearray.scala 134:13]
  wire  PENetwork_30_io_to_pes_1_out_valid; // @[pearray.scala 134:13]
  wire [7:0] PENetwork_30_io_to_pes_1_out_bits; // @[pearray.scala 134:13]
  wire  PENetwork_30_io_to_pes_2_in_valid; // @[pearray.scala 134:13]
  wire [7:0] PENetwork_30_io_to_pes_2_in_bits; // @[pearray.scala 134:13]
  wire  PENetwork_30_io_to_pes_2_out_valid; // @[pearray.scala 134:13]
  wire [7:0] PENetwork_30_io_to_pes_2_out_bits; // @[pearray.scala 134:13]
  wire  PENetwork_30_io_to_pes_3_in_valid; // @[pearray.scala 134:13]
  wire [7:0] PENetwork_30_io_to_pes_3_in_bits; // @[pearray.scala 134:13]
  wire  PENetwork_30_io_to_pes_3_out_valid; // @[pearray.scala 134:13]
  wire [7:0] PENetwork_30_io_to_pes_3_out_bits; // @[pearray.scala 134:13]
  wire  PENetwork_30_io_to_pes_4_in_valid; // @[pearray.scala 134:13]
  wire [7:0] PENetwork_30_io_to_pes_4_in_bits; // @[pearray.scala 134:13]
  wire  PENetwork_30_io_to_pes_4_out_valid; // @[pearray.scala 134:13]
  wire [7:0] PENetwork_30_io_to_pes_4_out_bits; // @[pearray.scala 134:13]
  wire  PENetwork_30_io_to_pes_5_in_valid; // @[pearray.scala 134:13]
  wire [7:0] PENetwork_30_io_to_pes_5_in_bits; // @[pearray.scala 134:13]
  wire  PENetwork_30_io_to_pes_5_out_valid; // @[pearray.scala 134:13]
  wire [7:0] PENetwork_30_io_to_pes_5_out_bits; // @[pearray.scala 134:13]
  wire  PENetwork_30_io_to_pes_6_in_valid; // @[pearray.scala 134:13]
  wire [7:0] PENetwork_30_io_to_pes_6_in_bits; // @[pearray.scala 134:13]
  wire  PENetwork_30_io_to_pes_6_out_valid; // @[pearray.scala 134:13]
  wire [7:0] PENetwork_30_io_to_pes_6_out_bits; // @[pearray.scala 134:13]
  wire  PENetwork_30_io_to_pes_7_in_valid; // @[pearray.scala 134:13]
  wire [7:0] PENetwork_30_io_to_pes_7_in_bits; // @[pearray.scala 134:13]
  wire  PENetwork_30_io_to_mem_valid; // @[pearray.scala 134:13]
  wire [7:0] PENetwork_30_io_to_mem_bits; // @[pearray.scala 134:13]
  wire  PENetwork_31_io_to_pes_0_in_valid; // @[pearray.scala 134:13]
  wire [7:0] PENetwork_31_io_to_pes_0_in_bits; // @[pearray.scala 134:13]
  wire  PENetwork_31_io_to_pes_0_out_valid; // @[pearray.scala 134:13]
  wire [7:0] PENetwork_31_io_to_pes_0_out_bits; // @[pearray.scala 134:13]
  wire  PENetwork_31_io_to_pes_1_in_valid; // @[pearray.scala 134:13]
  wire [7:0] PENetwork_31_io_to_pes_1_in_bits; // @[pearray.scala 134:13]
  wire  PENetwork_31_io_to_pes_1_out_valid; // @[pearray.scala 134:13]
  wire [7:0] PENetwork_31_io_to_pes_1_out_bits; // @[pearray.scala 134:13]
  wire  PENetwork_31_io_to_pes_2_in_valid; // @[pearray.scala 134:13]
  wire [7:0] PENetwork_31_io_to_pes_2_in_bits; // @[pearray.scala 134:13]
  wire  PENetwork_31_io_to_pes_2_out_valid; // @[pearray.scala 134:13]
  wire [7:0] PENetwork_31_io_to_pes_2_out_bits; // @[pearray.scala 134:13]
  wire  PENetwork_31_io_to_pes_3_in_valid; // @[pearray.scala 134:13]
  wire [7:0] PENetwork_31_io_to_pes_3_in_bits; // @[pearray.scala 134:13]
  wire  PENetwork_31_io_to_pes_3_out_valid; // @[pearray.scala 134:13]
  wire [7:0] PENetwork_31_io_to_pes_3_out_bits; // @[pearray.scala 134:13]
  wire  PENetwork_31_io_to_pes_4_in_valid; // @[pearray.scala 134:13]
  wire [7:0] PENetwork_31_io_to_pes_4_in_bits; // @[pearray.scala 134:13]
  wire  PENetwork_31_io_to_pes_4_out_valid; // @[pearray.scala 134:13]
  wire [7:0] PENetwork_31_io_to_pes_4_out_bits; // @[pearray.scala 134:13]
  wire  PENetwork_31_io_to_pes_5_in_valid; // @[pearray.scala 134:13]
  wire [7:0] PENetwork_31_io_to_pes_5_in_bits; // @[pearray.scala 134:13]
  wire  PENetwork_31_io_to_pes_5_out_valid; // @[pearray.scala 134:13]
  wire [7:0] PENetwork_31_io_to_pes_5_out_bits; // @[pearray.scala 134:13]
  wire  PENetwork_31_io_to_pes_6_in_valid; // @[pearray.scala 134:13]
  wire [7:0] PENetwork_31_io_to_pes_6_in_bits; // @[pearray.scala 134:13]
  wire  PENetwork_31_io_to_pes_6_out_valid; // @[pearray.scala 134:13]
  wire [7:0] PENetwork_31_io_to_pes_6_out_bits; // @[pearray.scala 134:13]
  wire  PENetwork_31_io_to_pes_7_in_valid; // @[pearray.scala 134:13]
  wire [7:0] PENetwork_31_io_to_pes_7_in_bits; // @[pearray.scala 134:13]
  wire  PENetwork_31_io_to_mem_valid; // @[pearray.scala 134:13]
  wire [7:0] PENetwork_31_io_to_mem_bits; // @[pearray.scala 134:13]
  wire [7:0] PENetwork_32_io_to_pes_0_in_bits; // @[pearray.scala 134:13]
  wire [7:0] PENetwork_32_io_to_pes_0_out_bits; // @[pearray.scala 134:13]
  wire [7:0] PENetwork_32_io_to_pes_1_in_bits; // @[pearray.scala 134:13]
  wire [7:0] PENetwork_32_io_to_pes_1_out_bits; // @[pearray.scala 134:13]
  wire [7:0] PENetwork_32_io_to_pes_2_in_bits; // @[pearray.scala 134:13]
  wire [7:0] PENetwork_32_io_to_pes_2_out_bits; // @[pearray.scala 134:13]
  wire [7:0] PENetwork_32_io_to_pes_3_in_bits; // @[pearray.scala 134:13]
  wire [7:0] PENetwork_32_io_to_pes_3_out_bits; // @[pearray.scala 134:13]
  wire [7:0] PENetwork_32_io_to_pes_4_in_bits; // @[pearray.scala 134:13]
  wire [7:0] PENetwork_32_io_to_pes_4_out_bits; // @[pearray.scala 134:13]
  wire [7:0] PENetwork_32_io_to_pes_5_in_bits; // @[pearray.scala 134:13]
  wire [7:0] PENetwork_32_io_to_pes_5_out_bits; // @[pearray.scala 134:13]
  wire [7:0] PENetwork_32_io_to_pes_6_in_bits; // @[pearray.scala 134:13]
  wire [7:0] PENetwork_32_io_to_pes_6_out_bits; // @[pearray.scala 134:13]
  wire [7:0] PENetwork_32_io_to_pes_7_in_bits; // @[pearray.scala 134:13]
  wire [7:0] PENetwork_32_io_to_pes_7_out_bits; // @[pearray.scala 134:13]
  wire [7:0] PENetwork_32_io_to_pes_8_in_bits; // @[pearray.scala 134:13]
  wire [7:0] PENetwork_32_io_to_pes_8_out_bits; // @[pearray.scala 134:13]
  wire [7:0] PENetwork_32_io_to_pes_9_in_bits; // @[pearray.scala 134:13]
  wire [7:0] PENetwork_32_io_to_pes_9_out_bits; // @[pearray.scala 134:13]
  wire [7:0] PENetwork_32_io_to_pes_10_in_bits; // @[pearray.scala 134:13]
  wire [7:0] PENetwork_32_io_to_pes_10_out_bits; // @[pearray.scala 134:13]
  wire [7:0] PENetwork_32_io_to_pes_11_in_bits; // @[pearray.scala 134:13]
  wire [7:0] PENetwork_32_io_to_pes_11_out_bits; // @[pearray.scala 134:13]
  wire [7:0] PENetwork_32_io_to_pes_12_in_bits; // @[pearray.scala 134:13]
  wire [7:0] PENetwork_32_io_to_pes_12_out_bits; // @[pearray.scala 134:13]
  wire [7:0] PENetwork_32_io_to_pes_13_in_bits; // @[pearray.scala 134:13]
  wire [7:0] PENetwork_32_io_to_pes_13_out_bits; // @[pearray.scala 134:13]
  wire [7:0] PENetwork_32_io_to_pes_14_in_bits; // @[pearray.scala 134:13]
  wire [7:0] PENetwork_32_io_to_pes_14_out_bits; // @[pearray.scala 134:13]
  wire [7:0] PENetwork_32_io_to_pes_15_in_bits; // @[pearray.scala 134:13]
  wire [7:0] PENetwork_32_io_to_mem_bits; // @[pearray.scala 134:13]
  wire [7:0] PENetwork_33_io_to_pes_0_in_bits; // @[pearray.scala 134:13]
  wire [7:0] PENetwork_33_io_to_pes_0_out_bits; // @[pearray.scala 134:13]
  wire [7:0] PENetwork_33_io_to_pes_1_in_bits; // @[pearray.scala 134:13]
  wire [7:0] PENetwork_33_io_to_pes_1_out_bits; // @[pearray.scala 134:13]
  wire [7:0] PENetwork_33_io_to_pes_2_in_bits; // @[pearray.scala 134:13]
  wire [7:0] PENetwork_33_io_to_pes_2_out_bits; // @[pearray.scala 134:13]
  wire [7:0] PENetwork_33_io_to_pes_3_in_bits; // @[pearray.scala 134:13]
  wire [7:0] PENetwork_33_io_to_pes_3_out_bits; // @[pearray.scala 134:13]
  wire [7:0] PENetwork_33_io_to_pes_4_in_bits; // @[pearray.scala 134:13]
  wire [7:0] PENetwork_33_io_to_pes_4_out_bits; // @[pearray.scala 134:13]
  wire [7:0] PENetwork_33_io_to_pes_5_in_bits; // @[pearray.scala 134:13]
  wire [7:0] PENetwork_33_io_to_pes_5_out_bits; // @[pearray.scala 134:13]
  wire [7:0] PENetwork_33_io_to_pes_6_in_bits; // @[pearray.scala 134:13]
  wire [7:0] PENetwork_33_io_to_pes_6_out_bits; // @[pearray.scala 134:13]
  wire [7:0] PENetwork_33_io_to_pes_7_in_bits; // @[pearray.scala 134:13]
  wire [7:0] PENetwork_33_io_to_pes_7_out_bits; // @[pearray.scala 134:13]
  wire [7:0] PENetwork_33_io_to_pes_8_in_bits; // @[pearray.scala 134:13]
  wire [7:0] PENetwork_33_io_to_pes_8_out_bits; // @[pearray.scala 134:13]
  wire [7:0] PENetwork_33_io_to_pes_9_in_bits; // @[pearray.scala 134:13]
  wire [7:0] PENetwork_33_io_to_pes_9_out_bits; // @[pearray.scala 134:13]
  wire [7:0] PENetwork_33_io_to_pes_10_in_bits; // @[pearray.scala 134:13]
  wire [7:0] PENetwork_33_io_to_pes_10_out_bits; // @[pearray.scala 134:13]
  wire [7:0] PENetwork_33_io_to_pes_11_in_bits; // @[pearray.scala 134:13]
  wire [7:0] PENetwork_33_io_to_pes_11_out_bits; // @[pearray.scala 134:13]
  wire [7:0] PENetwork_33_io_to_pes_12_in_bits; // @[pearray.scala 134:13]
  wire [7:0] PENetwork_33_io_to_pes_12_out_bits; // @[pearray.scala 134:13]
  wire [7:0] PENetwork_33_io_to_pes_13_in_bits; // @[pearray.scala 134:13]
  wire [7:0] PENetwork_33_io_to_pes_13_out_bits; // @[pearray.scala 134:13]
  wire [7:0] PENetwork_33_io_to_pes_14_in_bits; // @[pearray.scala 134:13]
  wire [7:0] PENetwork_33_io_to_pes_14_out_bits; // @[pearray.scala 134:13]
  wire [7:0] PENetwork_33_io_to_pes_15_in_bits; // @[pearray.scala 134:13]
  wire [7:0] PENetwork_33_io_to_mem_bits; // @[pearray.scala 134:13]
  wire [7:0] PENetwork_34_io_to_pes_0_in_bits; // @[pearray.scala 134:13]
  wire [7:0] PENetwork_34_io_to_pes_0_out_bits; // @[pearray.scala 134:13]
  wire [7:0] PENetwork_34_io_to_pes_1_in_bits; // @[pearray.scala 134:13]
  wire [7:0] PENetwork_34_io_to_pes_1_out_bits; // @[pearray.scala 134:13]
  wire [7:0] PENetwork_34_io_to_pes_2_in_bits; // @[pearray.scala 134:13]
  wire [7:0] PENetwork_34_io_to_pes_2_out_bits; // @[pearray.scala 134:13]
  wire [7:0] PENetwork_34_io_to_pes_3_in_bits; // @[pearray.scala 134:13]
  wire [7:0] PENetwork_34_io_to_pes_3_out_bits; // @[pearray.scala 134:13]
  wire [7:0] PENetwork_34_io_to_pes_4_in_bits; // @[pearray.scala 134:13]
  wire [7:0] PENetwork_34_io_to_pes_4_out_bits; // @[pearray.scala 134:13]
  wire [7:0] PENetwork_34_io_to_pes_5_in_bits; // @[pearray.scala 134:13]
  wire [7:0] PENetwork_34_io_to_pes_5_out_bits; // @[pearray.scala 134:13]
  wire [7:0] PENetwork_34_io_to_pes_6_in_bits; // @[pearray.scala 134:13]
  wire [7:0] PENetwork_34_io_to_pes_6_out_bits; // @[pearray.scala 134:13]
  wire [7:0] PENetwork_34_io_to_pes_7_in_bits; // @[pearray.scala 134:13]
  wire [7:0] PENetwork_34_io_to_pes_7_out_bits; // @[pearray.scala 134:13]
  wire [7:0] PENetwork_34_io_to_pes_8_in_bits; // @[pearray.scala 134:13]
  wire [7:0] PENetwork_34_io_to_pes_8_out_bits; // @[pearray.scala 134:13]
  wire [7:0] PENetwork_34_io_to_pes_9_in_bits; // @[pearray.scala 134:13]
  wire [7:0] PENetwork_34_io_to_pes_9_out_bits; // @[pearray.scala 134:13]
  wire [7:0] PENetwork_34_io_to_pes_10_in_bits; // @[pearray.scala 134:13]
  wire [7:0] PENetwork_34_io_to_pes_10_out_bits; // @[pearray.scala 134:13]
  wire [7:0] PENetwork_34_io_to_pes_11_in_bits; // @[pearray.scala 134:13]
  wire [7:0] PENetwork_34_io_to_pes_11_out_bits; // @[pearray.scala 134:13]
  wire [7:0] PENetwork_34_io_to_pes_12_in_bits; // @[pearray.scala 134:13]
  wire [7:0] PENetwork_34_io_to_pes_12_out_bits; // @[pearray.scala 134:13]
  wire [7:0] PENetwork_34_io_to_pes_13_in_bits; // @[pearray.scala 134:13]
  wire [7:0] PENetwork_34_io_to_pes_13_out_bits; // @[pearray.scala 134:13]
  wire [7:0] PENetwork_34_io_to_pes_14_in_bits; // @[pearray.scala 134:13]
  wire [7:0] PENetwork_34_io_to_pes_14_out_bits; // @[pearray.scala 134:13]
  wire [7:0] PENetwork_34_io_to_pes_15_in_bits; // @[pearray.scala 134:13]
  wire [7:0] PENetwork_34_io_to_mem_bits; // @[pearray.scala 134:13]
  wire [7:0] PENetwork_35_io_to_pes_0_in_bits; // @[pearray.scala 134:13]
  wire [7:0] PENetwork_35_io_to_pes_0_out_bits; // @[pearray.scala 134:13]
  wire [7:0] PENetwork_35_io_to_pes_1_in_bits; // @[pearray.scala 134:13]
  wire [7:0] PENetwork_35_io_to_pes_1_out_bits; // @[pearray.scala 134:13]
  wire [7:0] PENetwork_35_io_to_pes_2_in_bits; // @[pearray.scala 134:13]
  wire [7:0] PENetwork_35_io_to_pes_2_out_bits; // @[pearray.scala 134:13]
  wire [7:0] PENetwork_35_io_to_pes_3_in_bits; // @[pearray.scala 134:13]
  wire [7:0] PENetwork_35_io_to_pes_3_out_bits; // @[pearray.scala 134:13]
  wire [7:0] PENetwork_35_io_to_pes_4_in_bits; // @[pearray.scala 134:13]
  wire [7:0] PENetwork_35_io_to_pes_4_out_bits; // @[pearray.scala 134:13]
  wire [7:0] PENetwork_35_io_to_pes_5_in_bits; // @[pearray.scala 134:13]
  wire [7:0] PENetwork_35_io_to_pes_5_out_bits; // @[pearray.scala 134:13]
  wire [7:0] PENetwork_35_io_to_pes_6_in_bits; // @[pearray.scala 134:13]
  wire [7:0] PENetwork_35_io_to_pes_6_out_bits; // @[pearray.scala 134:13]
  wire [7:0] PENetwork_35_io_to_pes_7_in_bits; // @[pearray.scala 134:13]
  wire [7:0] PENetwork_35_io_to_pes_7_out_bits; // @[pearray.scala 134:13]
  wire [7:0] PENetwork_35_io_to_pes_8_in_bits; // @[pearray.scala 134:13]
  wire [7:0] PENetwork_35_io_to_pes_8_out_bits; // @[pearray.scala 134:13]
  wire [7:0] PENetwork_35_io_to_pes_9_in_bits; // @[pearray.scala 134:13]
  wire [7:0] PENetwork_35_io_to_pes_9_out_bits; // @[pearray.scala 134:13]
  wire [7:0] PENetwork_35_io_to_pes_10_in_bits; // @[pearray.scala 134:13]
  wire [7:0] PENetwork_35_io_to_pes_10_out_bits; // @[pearray.scala 134:13]
  wire [7:0] PENetwork_35_io_to_pes_11_in_bits; // @[pearray.scala 134:13]
  wire [7:0] PENetwork_35_io_to_pes_11_out_bits; // @[pearray.scala 134:13]
  wire [7:0] PENetwork_35_io_to_pes_12_in_bits; // @[pearray.scala 134:13]
  wire [7:0] PENetwork_35_io_to_pes_12_out_bits; // @[pearray.scala 134:13]
  wire [7:0] PENetwork_35_io_to_pes_13_in_bits; // @[pearray.scala 134:13]
  wire [7:0] PENetwork_35_io_to_pes_13_out_bits; // @[pearray.scala 134:13]
  wire [7:0] PENetwork_35_io_to_pes_14_in_bits; // @[pearray.scala 134:13]
  wire [7:0] PENetwork_35_io_to_pes_14_out_bits; // @[pearray.scala 134:13]
  wire [7:0] PENetwork_35_io_to_pes_15_in_bits; // @[pearray.scala 134:13]
  wire [7:0] PENetwork_35_io_to_mem_bits; // @[pearray.scala 134:13]
  wire [7:0] PENetwork_36_io_to_pes_0_in_bits; // @[pearray.scala 134:13]
  wire [7:0] PENetwork_36_io_to_pes_0_out_bits; // @[pearray.scala 134:13]
  wire [7:0] PENetwork_36_io_to_pes_1_in_bits; // @[pearray.scala 134:13]
  wire [7:0] PENetwork_36_io_to_pes_1_out_bits; // @[pearray.scala 134:13]
  wire [7:0] PENetwork_36_io_to_pes_2_in_bits; // @[pearray.scala 134:13]
  wire [7:0] PENetwork_36_io_to_pes_2_out_bits; // @[pearray.scala 134:13]
  wire [7:0] PENetwork_36_io_to_pes_3_in_bits; // @[pearray.scala 134:13]
  wire [7:0] PENetwork_36_io_to_pes_3_out_bits; // @[pearray.scala 134:13]
  wire [7:0] PENetwork_36_io_to_pes_4_in_bits; // @[pearray.scala 134:13]
  wire [7:0] PENetwork_36_io_to_pes_4_out_bits; // @[pearray.scala 134:13]
  wire [7:0] PENetwork_36_io_to_pes_5_in_bits; // @[pearray.scala 134:13]
  wire [7:0] PENetwork_36_io_to_pes_5_out_bits; // @[pearray.scala 134:13]
  wire [7:0] PENetwork_36_io_to_pes_6_in_bits; // @[pearray.scala 134:13]
  wire [7:0] PENetwork_36_io_to_pes_6_out_bits; // @[pearray.scala 134:13]
  wire [7:0] PENetwork_36_io_to_pes_7_in_bits; // @[pearray.scala 134:13]
  wire [7:0] PENetwork_36_io_to_pes_7_out_bits; // @[pearray.scala 134:13]
  wire [7:0] PENetwork_36_io_to_pes_8_in_bits; // @[pearray.scala 134:13]
  wire [7:0] PENetwork_36_io_to_pes_8_out_bits; // @[pearray.scala 134:13]
  wire [7:0] PENetwork_36_io_to_pes_9_in_bits; // @[pearray.scala 134:13]
  wire [7:0] PENetwork_36_io_to_pes_9_out_bits; // @[pearray.scala 134:13]
  wire [7:0] PENetwork_36_io_to_pes_10_in_bits; // @[pearray.scala 134:13]
  wire [7:0] PENetwork_36_io_to_pes_10_out_bits; // @[pearray.scala 134:13]
  wire [7:0] PENetwork_36_io_to_pes_11_in_bits; // @[pearray.scala 134:13]
  wire [7:0] PENetwork_36_io_to_pes_11_out_bits; // @[pearray.scala 134:13]
  wire [7:0] PENetwork_36_io_to_pes_12_in_bits; // @[pearray.scala 134:13]
  wire [7:0] PENetwork_36_io_to_pes_12_out_bits; // @[pearray.scala 134:13]
  wire [7:0] PENetwork_36_io_to_pes_13_in_bits; // @[pearray.scala 134:13]
  wire [7:0] PENetwork_36_io_to_pes_13_out_bits; // @[pearray.scala 134:13]
  wire [7:0] PENetwork_36_io_to_pes_14_in_bits; // @[pearray.scala 134:13]
  wire [7:0] PENetwork_36_io_to_pes_14_out_bits; // @[pearray.scala 134:13]
  wire [7:0] PENetwork_36_io_to_pes_15_in_bits; // @[pearray.scala 134:13]
  wire [7:0] PENetwork_36_io_to_mem_bits; // @[pearray.scala 134:13]
  wire [7:0] PENetwork_37_io_to_pes_0_in_bits; // @[pearray.scala 134:13]
  wire [7:0] PENetwork_37_io_to_pes_0_out_bits; // @[pearray.scala 134:13]
  wire [7:0] PENetwork_37_io_to_pes_1_in_bits; // @[pearray.scala 134:13]
  wire [7:0] PENetwork_37_io_to_pes_1_out_bits; // @[pearray.scala 134:13]
  wire [7:0] PENetwork_37_io_to_pes_2_in_bits; // @[pearray.scala 134:13]
  wire [7:0] PENetwork_37_io_to_pes_2_out_bits; // @[pearray.scala 134:13]
  wire [7:0] PENetwork_37_io_to_pes_3_in_bits; // @[pearray.scala 134:13]
  wire [7:0] PENetwork_37_io_to_pes_3_out_bits; // @[pearray.scala 134:13]
  wire [7:0] PENetwork_37_io_to_pes_4_in_bits; // @[pearray.scala 134:13]
  wire [7:0] PENetwork_37_io_to_pes_4_out_bits; // @[pearray.scala 134:13]
  wire [7:0] PENetwork_37_io_to_pes_5_in_bits; // @[pearray.scala 134:13]
  wire [7:0] PENetwork_37_io_to_pes_5_out_bits; // @[pearray.scala 134:13]
  wire [7:0] PENetwork_37_io_to_pes_6_in_bits; // @[pearray.scala 134:13]
  wire [7:0] PENetwork_37_io_to_pes_6_out_bits; // @[pearray.scala 134:13]
  wire [7:0] PENetwork_37_io_to_pes_7_in_bits; // @[pearray.scala 134:13]
  wire [7:0] PENetwork_37_io_to_pes_7_out_bits; // @[pearray.scala 134:13]
  wire [7:0] PENetwork_37_io_to_pes_8_in_bits; // @[pearray.scala 134:13]
  wire [7:0] PENetwork_37_io_to_pes_8_out_bits; // @[pearray.scala 134:13]
  wire [7:0] PENetwork_37_io_to_pes_9_in_bits; // @[pearray.scala 134:13]
  wire [7:0] PENetwork_37_io_to_pes_9_out_bits; // @[pearray.scala 134:13]
  wire [7:0] PENetwork_37_io_to_pes_10_in_bits; // @[pearray.scala 134:13]
  wire [7:0] PENetwork_37_io_to_pes_10_out_bits; // @[pearray.scala 134:13]
  wire [7:0] PENetwork_37_io_to_pes_11_in_bits; // @[pearray.scala 134:13]
  wire [7:0] PENetwork_37_io_to_pes_11_out_bits; // @[pearray.scala 134:13]
  wire [7:0] PENetwork_37_io_to_pes_12_in_bits; // @[pearray.scala 134:13]
  wire [7:0] PENetwork_37_io_to_pes_12_out_bits; // @[pearray.scala 134:13]
  wire [7:0] PENetwork_37_io_to_pes_13_in_bits; // @[pearray.scala 134:13]
  wire [7:0] PENetwork_37_io_to_pes_13_out_bits; // @[pearray.scala 134:13]
  wire [7:0] PENetwork_37_io_to_pes_14_in_bits; // @[pearray.scala 134:13]
  wire [7:0] PENetwork_37_io_to_pes_14_out_bits; // @[pearray.scala 134:13]
  wire [7:0] PENetwork_37_io_to_pes_15_in_bits; // @[pearray.scala 134:13]
  wire [7:0] PENetwork_37_io_to_mem_bits; // @[pearray.scala 134:13]
  wire [7:0] PENetwork_38_io_to_pes_0_in_bits; // @[pearray.scala 134:13]
  wire [7:0] PENetwork_38_io_to_pes_0_out_bits; // @[pearray.scala 134:13]
  wire [7:0] PENetwork_38_io_to_pes_1_in_bits; // @[pearray.scala 134:13]
  wire [7:0] PENetwork_38_io_to_pes_1_out_bits; // @[pearray.scala 134:13]
  wire [7:0] PENetwork_38_io_to_pes_2_in_bits; // @[pearray.scala 134:13]
  wire [7:0] PENetwork_38_io_to_pes_2_out_bits; // @[pearray.scala 134:13]
  wire [7:0] PENetwork_38_io_to_pes_3_in_bits; // @[pearray.scala 134:13]
  wire [7:0] PENetwork_38_io_to_pes_3_out_bits; // @[pearray.scala 134:13]
  wire [7:0] PENetwork_38_io_to_pes_4_in_bits; // @[pearray.scala 134:13]
  wire [7:0] PENetwork_38_io_to_pes_4_out_bits; // @[pearray.scala 134:13]
  wire [7:0] PENetwork_38_io_to_pes_5_in_bits; // @[pearray.scala 134:13]
  wire [7:0] PENetwork_38_io_to_pes_5_out_bits; // @[pearray.scala 134:13]
  wire [7:0] PENetwork_38_io_to_pes_6_in_bits; // @[pearray.scala 134:13]
  wire [7:0] PENetwork_38_io_to_pes_6_out_bits; // @[pearray.scala 134:13]
  wire [7:0] PENetwork_38_io_to_pes_7_in_bits; // @[pearray.scala 134:13]
  wire [7:0] PENetwork_38_io_to_pes_7_out_bits; // @[pearray.scala 134:13]
  wire [7:0] PENetwork_38_io_to_pes_8_in_bits; // @[pearray.scala 134:13]
  wire [7:0] PENetwork_38_io_to_pes_8_out_bits; // @[pearray.scala 134:13]
  wire [7:0] PENetwork_38_io_to_pes_9_in_bits; // @[pearray.scala 134:13]
  wire [7:0] PENetwork_38_io_to_pes_9_out_bits; // @[pearray.scala 134:13]
  wire [7:0] PENetwork_38_io_to_pes_10_in_bits; // @[pearray.scala 134:13]
  wire [7:0] PENetwork_38_io_to_pes_10_out_bits; // @[pearray.scala 134:13]
  wire [7:0] PENetwork_38_io_to_pes_11_in_bits; // @[pearray.scala 134:13]
  wire [7:0] PENetwork_38_io_to_pes_11_out_bits; // @[pearray.scala 134:13]
  wire [7:0] PENetwork_38_io_to_pes_12_in_bits; // @[pearray.scala 134:13]
  wire [7:0] PENetwork_38_io_to_pes_12_out_bits; // @[pearray.scala 134:13]
  wire [7:0] PENetwork_38_io_to_pes_13_in_bits; // @[pearray.scala 134:13]
  wire [7:0] PENetwork_38_io_to_pes_13_out_bits; // @[pearray.scala 134:13]
  wire [7:0] PENetwork_38_io_to_pes_14_in_bits; // @[pearray.scala 134:13]
  wire [7:0] PENetwork_38_io_to_pes_14_out_bits; // @[pearray.scala 134:13]
  wire [7:0] PENetwork_38_io_to_pes_15_in_bits; // @[pearray.scala 134:13]
  wire [7:0] PENetwork_38_io_to_mem_bits; // @[pearray.scala 134:13]
  wire [7:0] PENetwork_39_io_to_pes_0_in_bits; // @[pearray.scala 134:13]
  wire [7:0] PENetwork_39_io_to_pes_0_out_bits; // @[pearray.scala 134:13]
  wire [7:0] PENetwork_39_io_to_pes_1_in_bits; // @[pearray.scala 134:13]
  wire [7:0] PENetwork_39_io_to_pes_1_out_bits; // @[pearray.scala 134:13]
  wire [7:0] PENetwork_39_io_to_pes_2_in_bits; // @[pearray.scala 134:13]
  wire [7:0] PENetwork_39_io_to_pes_2_out_bits; // @[pearray.scala 134:13]
  wire [7:0] PENetwork_39_io_to_pes_3_in_bits; // @[pearray.scala 134:13]
  wire [7:0] PENetwork_39_io_to_pes_3_out_bits; // @[pearray.scala 134:13]
  wire [7:0] PENetwork_39_io_to_pes_4_in_bits; // @[pearray.scala 134:13]
  wire [7:0] PENetwork_39_io_to_pes_4_out_bits; // @[pearray.scala 134:13]
  wire [7:0] PENetwork_39_io_to_pes_5_in_bits; // @[pearray.scala 134:13]
  wire [7:0] PENetwork_39_io_to_pes_5_out_bits; // @[pearray.scala 134:13]
  wire [7:0] PENetwork_39_io_to_pes_6_in_bits; // @[pearray.scala 134:13]
  wire [7:0] PENetwork_39_io_to_pes_6_out_bits; // @[pearray.scala 134:13]
  wire [7:0] PENetwork_39_io_to_pes_7_in_bits; // @[pearray.scala 134:13]
  wire [7:0] PENetwork_39_io_to_pes_7_out_bits; // @[pearray.scala 134:13]
  wire [7:0] PENetwork_39_io_to_pes_8_in_bits; // @[pearray.scala 134:13]
  wire [7:0] PENetwork_39_io_to_pes_8_out_bits; // @[pearray.scala 134:13]
  wire [7:0] PENetwork_39_io_to_pes_9_in_bits; // @[pearray.scala 134:13]
  wire [7:0] PENetwork_39_io_to_pes_9_out_bits; // @[pearray.scala 134:13]
  wire [7:0] PENetwork_39_io_to_pes_10_in_bits; // @[pearray.scala 134:13]
  wire [7:0] PENetwork_39_io_to_pes_10_out_bits; // @[pearray.scala 134:13]
  wire [7:0] PENetwork_39_io_to_pes_11_in_bits; // @[pearray.scala 134:13]
  wire [7:0] PENetwork_39_io_to_pes_11_out_bits; // @[pearray.scala 134:13]
  wire [7:0] PENetwork_39_io_to_pes_12_in_bits; // @[pearray.scala 134:13]
  wire [7:0] PENetwork_39_io_to_pes_12_out_bits; // @[pearray.scala 134:13]
  wire [7:0] PENetwork_39_io_to_pes_13_in_bits; // @[pearray.scala 134:13]
  wire [7:0] PENetwork_39_io_to_pes_13_out_bits; // @[pearray.scala 134:13]
  wire [7:0] PENetwork_39_io_to_pes_14_in_bits; // @[pearray.scala 134:13]
  wire [7:0] PENetwork_39_io_to_pes_14_out_bits; // @[pearray.scala 134:13]
  wire [7:0] PENetwork_39_io_to_pes_15_in_bits; // @[pearray.scala 134:13]
  wire [7:0] PENetwork_39_io_to_mem_bits; // @[pearray.scala 134:13]
  wire  MemController_clock; // @[pearray.scala 202:15]
  wire  MemController_reset; // @[pearray.scala 202:15]
  wire  MemController_io_rd_valid; // @[pearray.scala 202:15]
  wire  MemController_io_wr_valid; // @[pearray.scala 202:15]
  wire  MemController_io_rd_data_valid; // @[pearray.scala 202:15]
  wire [7:0] MemController_io_rd_data_bits; // @[pearray.scala 202:15]
  wire  MemController_io_wr_data_valid; // @[pearray.scala 202:15]
  wire [7:0] MemController_io_wr_data_bits; // @[pearray.scala 202:15]
  wire  MemController_1_clock; // @[pearray.scala 202:15]
  wire  MemController_1_reset; // @[pearray.scala 202:15]
  wire  MemController_1_io_rd_valid; // @[pearray.scala 202:15]
  wire  MemController_1_io_wr_valid; // @[pearray.scala 202:15]
  wire  MemController_1_io_rd_data_valid; // @[pearray.scala 202:15]
  wire [7:0] MemController_1_io_rd_data_bits; // @[pearray.scala 202:15]
  wire  MemController_1_io_wr_data_valid; // @[pearray.scala 202:15]
  wire [7:0] MemController_1_io_wr_data_bits; // @[pearray.scala 202:15]
  wire  MemController_2_clock; // @[pearray.scala 202:15]
  wire  MemController_2_reset; // @[pearray.scala 202:15]
  wire  MemController_2_io_rd_valid; // @[pearray.scala 202:15]
  wire  MemController_2_io_wr_valid; // @[pearray.scala 202:15]
  wire  MemController_2_io_rd_data_valid; // @[pearray.scala 202:15]
  wire [7:0] MemController_2_io_rd_data_bits; // @[pearray.scala 202:15]
  wire  MemController_2_io_wr_data_valid; // @[pearray.scala 202:15]
  wire [7:0] MemController_2_io_wr_data_bits; // @[pearray.scala 202:15]
  wire  MemController_3_clock; // @[pearray.scala 202:15]
  wire  MemController_3_reset; // @[pearray.scala 202:15]
  wire  MemController_3_io_rd_valid; // @[pearray.scala 202:15]
  wire  MemController_3_io_wr_valid; // @[pearray.scala 202:15]
  wire  MemController_3_io_rd_data_valid; // @[pearray.scala 202:15]
  wire [7:0] MemController_3_io_rd_data_bits; // @[pearray.scala 202:15]
  wire  MemController_3_io_wr_data_valid; // @[pearray.scala 202:15]
  wire [7:0] MemController_3_io_wr_data_bits; // @[pearray.scala 202:15]
  wire  MemController_4_clock; // @[pearray.scala 202:15]
  wire  MemController_4_reset; // @[pearray.scala 202:15]
  wire  MemController_4_io_rd_valid; // @[pearray.scala 202:15]
  wire  MemController_4_io_wr_valid; // @[pearray.scala 202:15]
  wire  MemController_4_io_rd_data_valid; // @[pearray.scala 202:15]
  wire [7:0] MemController_4_io_rd_data_bits; // @[pearray.scala 202:15]
  wire  MemController_4_io_wr_data_valid; // @[pearray.scala 202:15]
  wire [7:0] MemController_4_io_wr_data_bits; // @[pearray.scala 202:15]
  wire  MemController_5_clock; // @[pearray.scala 202:15]
  wire  MemController_5_reset; // @[pearray.scala 202:15]
  wire  MemController_5_io_rd_valid; // @[pearray.scala 202:15]
  wire  MemController_5_io_wr_valid; // @[pearray.scala 202:15]
  wire  MemController_5_io_rd_data_valid; // @[pearray.scala 202:15]
  wire [7:0] MemController_5_io_rd_data_bits; // @[pearray.scala 202:15]
  wire  MemController_5_io_wr_data_valid; // @[pearray.scala 202:15]
  wire [7:0] MemController_5_io_wr_data_bits; // @[pearray.scala 202:15]
  wire  MemController_6_clock; // @[pearray.scala 202:15]
  wire  MemController_6_reset; // @[pearray.scala 202:15]
  wire  MemController_6_io_rd_valid; // @[pearray.scala 202:15]
  wire  MemController_6_io_wr_valid; // @[pearray.scala 202:15]
  wire  MemController_6_io_rd_data_valid; // @[pearray.scala 202:15]
  wire [7:0] MemController_6_io_rd_data_bits; // @[pearray.scala 202:15]
  wire  MemController_6_io_wr_data_valid; // @[pearray.scala 202:15]
  wire [7:0] MemController_6_io_wr_data_bits; // @[pearray.scala 202:15]
  wire  MemController_7_clock; // @[pearray.scala 202:15]
  wire  MemController_7_reset; // @[pearray.scala 202:15]
  wire  MemController_7_io_rd_valid; // @[pearray.scala 202:15]
  wire  MemController_7_io_wr_valid; // @[pearray.scala 202:15]
  wire  MemController_7_io_rd_data_valid; // @[pearray.scala 202:15]
  wire [7:0] MemController_7_io_rd_data_bits; // @[pearray.scala 202:15]
  wire  MemController_7_io_wr_data_valid; // @[pearray.scala 202:15]
  wire [7:0] MemController_7_io_wr_data_bits; // @[pearray.scala 202:15]
  wire  MemController_8_clock; // @[pearray.scala 202:15]
  wire  MemController_8_reset; // @[pearray.scala 202:15]
  wire  MemController_8_io_rd_valid; // @[pearray.scala 202:15]
  wire  MemController_8_io_wr_valid; // @[pearray.scala 202:15]
  wire  MemController_8_io_rd_data_valid; // @[pearray.scala 202:15]
  wire [7:0] MemController_8_io_rd_data_bits; // @[pearray.scala 202:15]
  wire  MemController_8_io_wr_data_valid; // @[pearray.scala 202:15]
  wire [7:0] MemController_8_io_wr_data_bits; // @[pearray.scala 202:15]
  wire  MemController_9_clock; // @[pearray.scala 202:15]
  wire  MemController_9_reset; // @[pearray.scala 202:15]
  wire  MemController_9_io_rd_valid; // @[pearray.scala 202:15]
  wire  MemController_9_io_wr_valid; // @[pearray.scala 202:15]
  wire  MemController_9_io_rd_data_valid; // @[pearray.scala 202:15]
  wire [7:0] MemController_9_io_rd_data_bits; // @[pearray.scala 202:15]
  wire  MemController_9_io_wr_data_valid; // @[pearray.scala 202:15]
  wire [7:0] MemController_9_io_wr_data_bits; // @[pearray.scala 202:15]
  wire  MemController_10_clock; // @[pearray.scala 202:15]
  wire  MemController_10_reset; // @[pearray.scala 202:15]
  wire  MemController_10_io_rd_valid; // @[pearray.scala 202:15]
  wire  MemController_10_io_wr_valid; // @[pearray.scala 202:15]
  wire  MemController_10_io_rd_data_valid; // @[pearray.scala 202:15]
  wire [7:0] MemController_10_io_rd_data_bits; // @[pearray.scala 202:15]
  wire  MemController_10_io_wr_data_valid; // @[pearray.scala 202:15]
  wire [7:0] MemController_10_io_wr_data_bits; // @[pearray.scala 202:15]
  wire  MemController_11_clock; // @[pearray.scala 202:15]
  wire  MemController_11_reset; // @[pearray.scala 202:15]
  wire  MemController_11_io_rd_valid; // @[pearray.scala 202:15]
  wire  MemController_11_io_wr_valid; // @[pearray.scala 202:15]
  wire  MemController_11_io_rd_data_valid; // @[pearray.scala 202:15]
  wire [7:0] MemController_11_io_rd_data_bits; // @[pearray.scala 202:15]
  wire  MemController_11_io_wr_data_valid; // @[pearray.scala 202:15]
  wire [7:0] MemController_11_io_wr_data_bits; // @[pearray.scala 202:15]
  wire  MemController_12_clock; // @[pearray.scala 202:15]
  wire  MemController_12_reset; // @[pearray.scala 202:15]
  wire  MemController_12_io_rd_valid; // @[pearray.scala 202:15]
  wire  MemController_12_io_wr_valid; // @[pearray.scala 202:15]
  wire  MemController_12_io_rd_data_valid; // @[pearray.scala 202:15]
  wire [7:0] MemController_12_io_rd_data_bits; // @[pearray.scala 202:15]
  wire  MemController_12_io_wr_data_valid; // @[pearray.scala 202:15]
  wire [7:0] MemController_12_io_wr_data_bits; // @[pearray.scala 202:15]
  wire  MemController_13_clock; // @[pearray.scala 202:15]
  wire  MemController_13_reset; // @[pearray.scala 202:15]
  wire  MemController_13_io_rd_valid; // @[pearray.scala 202:15]
  wire  MemController_13_io_wr_valid; // @[pearray.scala 202:15]
  wire  MemController_13_io_rd_data_valid; // @[pearray.scala 202:15]
  wire [7:0] MemController_13_io_rd_data_bits; // @[pearray.scala 202:15]
  wire  MemController_13_io_wr_data_valid; // @[pearray.scala 202:15]
  wire [7:0] MemController_13_io_wr_data_bits; // @[pearray.scala 202:15]
  wire  MemController_14_clock; // @[pearray.scala 202:15]
  wire  MemController_14_reset; // @[pearray.scala 202:15]
  wire  MemController_14_io_rd_valid; // @[pearray.scala 202:15]
  wire  MemController_14_io_wr_valid; // @[pearray.scala 202:15]
  wire  MemController_14_io_rd_data_valid; // @[pearray.scala 202:15]
  wire [7:0] MemController_14_io_rd_data_bits; // @[pearray.scala 202:15]
  wire  MemController_14_io_wr_data_valid; // @[pearray.scala 202:15]
  wire [7:0] MemController_14_io_wr_data_bits; // @[pearray.scala 202:15]
  wire  MemController_15_clock; // @[pearray.scala 202:15]
  wire  MemController_15_reset; // @[pearray.scala 202:15]
  wire  MemController_15_io_rd_valid; // @[pearray.scala 202:15]
  wire  MemController_15_io_wr_valid; // @[pearray.scala 202:15]
  wire  MemController_15_io_rd_data_valid; // @[pearray.scala 202:15]
  wire [7:0] MemController_15_io_rd_data_bits; // @[pearray.scala 202:15]
  wire  MemController_15_io_wr_data_valid; // @[pearray.scala 202:15]
  wire [7:0] MemController_15_io_wr_data_bits; // @[pearray.scala 202:15]
  wire  MemController_16_clock; // @[pearray.scala 200:15]
  wire  MemController_16_reset; // @[pearray.scala 200:15]
  wire  MemController_16_io_rd_valid; // @[pearray.scala 200:15]
  wire  MemController_16_io_wr_valid; // @[pearray.scala 200:15]
  wire  MemController_16_io_rd_data_valid; // @[pearray.scala 200:15]
  wire [7:0] MemController_16_io_rd_data_bits; // @[pearray.scala 200:15]
  wire  MemController_16_io_wr_data_valid; // @[pearray.scala 200:15]
  wire [7:0] MemController_16_io_wr_data_bits; // @[pearray.scala 200:15]
  wire  MemController_17_clock; // @[pearray.scala 200:15]
  wire  MemController_17_reset; // @[pearray.scala 200:15]
  wire  MemController_17_io_rd_valid; // @[pearray.scala 200:15]
  wire  MemController_17_io_wr_valid; // @[pearray.scala 200:15]
  wire  MemController_17_io_rd_data_valid; // @[pearray.scala 200:15]
  wire [7:0] MemController_17_io_rd_data_bits; // @[pearray.scala 200:15]
  wire  MemController_17_io_wr_data_valid; // @[pearray.scala 200:15]
  wire [7:0] MemController_17_io_wr_data_bits; // @[pearray.scala 200:15]
  wire  MemController_18_clock; // @[pearray.scala 200:15]
  wire  MemController_18_reset; // @[pearray.scala 200:15]
  wire  MemController_18_io_rd_valid; // @[pearray.scala 200:15]
  wire  MemController_18_io_wr_valid; // @[pearray.scala 200:15]
  wire  MemController_18_io_rd_data_valid; // @[pearray.scala 200:15]
  wire [7:0] MemController_18_io_rd_data_bits; // @[pearray.scala 200:15]
  wire  MemController_18_io_wr_data_valid; // @[pearray.scala 200:15]
  wire [7:0] MemController_18_io_wr_data_bits; // @[pearray.scala 200:15]
  wire  MemController_19_clock; // @[pearray.scala 200:15]
  wire  MemController_19_reset; // @[pearray.scala 200:15]
  wire  MemController_19_io_rd_valid; // @[pearray.scala 200:15]
  wire  MemController_19_io_wr_valid; // @[pearray.scala 200:15]
  wire  MemController_19_io_rd_data_valid; // @[pearray.scala 200:15]
  wire [7:0] MemController_19_io_rd_data_bits; // @[pearray.scala 200:15]
  wire  MemController_19_io_wr_data_valid; // @[pearray.scala 200:15]
  wire [7:0] MemController_19_io_wr_data_bits; // @[pearray.scala 200:15]
  wire  MemController_20_clock; // @[pearray.scala 200:15]
  wire  MemController_20_reset; // @[pearray.scala 200:15]
  wire  MemController_20_io_rd_valid; // @[pearray.scala 200:15]
  wire  MemController_20_io_wr_valid; // @[pearray.scala 200:15]
  wire  MemController_20_io_rd_data_valid; // @[pearray.scala 200:15]
  wire [7:0] MemController_20_io_rd_data_bits; // @[pearray.scala 200:15]
  wire  MemController_20_io_wr_data_valid; // @[pearray.scala 200:15]
  wire [7:0] MemController_20_io_wr_data_bits; // @[pearray.scala 200:15]
  wire  MemController_21_clock; // @[pearray.scala 200:15]
  wire  MemController_21_reset; // @[pearray.scala 200:15]
  wire  MemController_21_io_rd_valid; // @[pearray.scala 200:15]
  wire  MemController_21_io_wr_valid; // @[pearray.scala 200:15]
  wire  MemController_21_io_rd_data_valid; // @[pearray.scala 200:15]
  wire [7:0] MemController_21_io_rd_data_bits; // @[pearray.scala 200:15]
  wire  MemController_21_io_wr_data_valid; // @[pearray.scala 200:15]
  wire [7:0] MemController_21_io_wr_data_bits; // @[pearray.scala 200:15]
  wire  MemController_22_clock; // @[pearray.scala 200:15]
  wire  MemController_22_reset; // @[pearray.scala 200:15]
  wire  MemController_22_io_rd_valid; // @[pearray.scala 200:15]
  wire  MemController_22_io_wr_valid; // @[pearray.scala 200:15]
  wire  MemController_22_io_rd_data_valid; // @[pearray.scala 200:15]
  wire [7:0] MemController_22_io_rd_data_bits; // @[pearray.scala 200:15]
  wire  MemController_22_io_wr_data_valid; // @[pearray.scala 200:15]
  wire [7:0] MemController_22_io_wr_data_bits; // @[pearray.scala 200:15]
  wire  MemController_23_clock; // @[pearray.scala 200:15]
  wire  MemController_23_reset; // @[pearray.scala 200:15]
  wire  MemController_23_io_rd_valid; // @[pearray.scala 200:15]
  wire  MemController_23_io_wr_valid; // @[pearray.scala 200:15]
  wire  MemController_23_io_rd_data_valid; // @[pearray.scala 200:15]
  wire [7:0] MemController_23_io_rd_data_bits; // @[pearray.scala 200:15]
  wire  MemController_23_io_wr_data_valid; // @[pearray.scala 200:15]
  wire [7:0] MemController_23_io_wr_data_bits; // @[pearray.scala 200:15]
  wire  MemController_24_clock; // @[pearray.scala 200:15]
  wire  MemController_24_reset; // @[pearray.scala 200:15]
  wire  MemController_24_io_rd_valid; // @[pearray.scala 200:15]
  wire  MemController_24_io_wr_valid; // @[pearray.scala 200:15]
  wire  MemController_24_io_rd_data_valid; // @[pearray.scala 200:15]
  wire [7:0] MemController_24_io_rd_data_bits; // @[pearray.scala 200:15]
  wire  MemController_24_io_wr_data_valid; // @[pearray.scala 200:15]
  wire [7:0] MemController_24_io_wr_data_bits; // @[pearray.scala 200:15]
  wire  MemController_25_clock; // @[pearray.scala 200:15]
  wire  MemController_25_reset; // @[pearray.scala 200:15]
  wire  MemController_25_io_rd_valid; // @[pearray.scala 200:15]
  wire  MemController_25_io_wr_valid; // @[pearray.scala 200:15]
  wire  MemController_25_io_rd_data_valid; // @[pearray.scala 200:15]
  wire [7:0] MemController_25_io_rd_data_bits; // @[pearray.scala 200:15]
  wire  MemController_25_io_wr_data_valid; // @[pearray.scala 200:15]
  wire [7:0] MemController_25_io_wr_data_bits; // @[pearray.scala 200:15]
  wire  MemController_26_clock; // @[pearray.scala 200:15]
  wire  MemController_26_reset; // @[pearray.scala 200:15]
  wire  MemController_26_io_rd_valid; // @[pearray.scala 200:15]
  wire  MemController_26_io_wr_valid; // @[pearray.scala 200:15]
  wire  MemController_26_io_rd_data_valid; // @[pearray.scala 200:15]
  wire [7:0] MemController_26_io_rd_data_bits; // @[pearray.scala 200:15]
  wire  MemController_26_io_wr_data_valid; // @[pearray.scala 200:15]
  wire [7:0] MemController_26_io_wr_data_bits; // @[pearray.scala 200:15]
  wire  MemController_27_clock; // @[pearray.scala 200:15]
  wire  MemController_27_reset; // @[pearray.scala 200:15]
  wire  MemController_27_io_rd_valid; // @[pearray.scala 200:15]
  wire  MemController_27_io_wr_valid; // @[pearray.scala 200:15]
  wire  MemController_27_io_rd_data_valid; // @[pearray.scala 200:15]
  wire [7:0] MemController_27_io_rd_data_bits; // @[pearray.scala 200:15]
  wire  MemController_27_io_wr_data_valid; // @[pearray.scala 200:15]
  wire [7:0] MemController_27_io_wr_data_bits; // @[pearray.scala 200:15]
  wire  MemController_28_clock; // @[pearray.scala 200:15]
  wire  MemController_28_reset; // @[pearray.scala 200:15]
  wire  MemController_28_io_rd_valid; // @[pearray.scala 200:15]
  wire  MemController_28_io_wr_valid; // @[pearray.scala 200:15]
  wire  MemController_28_io_rd_data_valid; // @[pearray.scala 200:15]
  wire [7:0] MemController_28_io_rd_data_bits; // @[pearray.scala 200:15]
  wire  MemController_28_io_wr_data_valid; // @[pearray.scala 200:15]
  wire [7:0] MemController_28_io_wr_data_bits; // @[pearray.scala 200:15]
  wire  MemController_29_clock; // @[pearray.scala 200:15]
  wire  MemController_29_reset; // @[pearray.scala 200:15]
  wire  MemController_29_io_rd_valid; // @[pearray.scala 200:15]
  wire  MemController_29_io_wr_valid; // @[pearray.scala 200:15]
  wire  MemController_29_io_rd_data_valid; // @[pearray.scala 200:15]
  wire [7:0] MemController_29_io_rd_data_bits; // @[pearray.scala 200:15]
  wire  MemController_29_io_wr_data_valid; // @[pearray.scala 200:15]
  wire [7:0] MemController_29_io_wr_data_bits; // @[pearray.scala 200:15]
  wire  MemController_30_clock; // @[pearray.scala 200:15]
  wire  MemController_30_reset; // @[pearray.scala 200:15]
  wire  MemController_30_io_rd_valid; // @[pearray.scala 200:15]
  wire  MemController_30_io_wr_valid; // @[pearray.scala 200:15]
  wire  MemController_30_io_rd_data_valid; // @[pearray.scala 200:15]
  wire [7:0] MemController_30_io_rd_data_bits; // @[pearray.scala 200:15]
  wire  MemController_30_io_wr_data_valid; // @[pearray.scala 200:15]
  wire [7:0] MemController_30_io_wr_data_bits; // @[pearray.scala 200:15]
  wire  MemController_31_clock; // @[pearray.scala 200:15]
  wire  MemController_31_reset; // @[pearray.scala 200:15]
  wire  MemController_31_io_rd_valid; // @[pearray.scala 200:15]
  wire  MemController_31_io_wr_valid; // @[pearray.scala 200:15]
  wire  MemController_31_io_rd_data_valid; // @[pearray.scala 200:15]
  wire [7:0] MemController_31_io_rd_data_bits; // @[pearray.scala 200:15]
  wire  MemController_31_io_wr_data_valid; // @[pearray.scala 200:15]
  wire [7:0] MemController_31_io_wr_data_bits; // @[pearray.scala 200:15]
  wire  MemController_32_clock; // @[pearray.scala 200:15]
  wire  MemController_32_reset; // @[pearray.scala 200:15]
  wire  MemController_32_io_rd_valid; // @[pearray.scala 200:15]
  wire  MemController_32_io_wr_valid; // @[pearray.scala 200:15]
  wire  MemController_32_io_rd_data_valid; // @[pearray.scala 200:15]
  wire [7:0] MemController_32_io_rd_data_bits; // @[pearray.scala 200:15]
  wire  MemController_32_io_wr_data_valid; // @[pearray.scala 200:15]
  wire [7:0] MemController_32_io_wr_data_bits; // @[pearray.scala 200:15]
  wire  MemController_33_clock; // @[pearray.scala 200:15]
  wire  MemController_33_reset; // @[pearray.scala 200:15]
  wire  MemController_33_io_rd_valid; // @[pearray.scala 200:15]
  wire  MemController_33_io_wr_valid; // @[pearray.scala 200:15]
  wire  MemController_33_io_rd_data_valid; // @[pearray.scala 200:15]
  wire [7:0] MemController_33_io_rd_data_bits; // @[pearray.scala 200:15]
  wire  MemController_33_io_wr_data_valid; // @[pearray.scala 200:15]
  wire [7:0] MemController_33_io_wr_data_bits; // @[pearray.scala 200:15]
  wire  MemController_34_clock; // @[pearray.scala 200:15]
  wire  MemController_34_reset; // @[pearray.scala 200:15]
  wire  MemController_34_io_rd_valid; // @[pearray.scala 200:15]
  wire  MemController_34_io_wr_valid; // @[pearray.scala 200:15]
  wire  MemController_34_io_rd_data_valid; // @[pearray.scala 200:15]
  wire [7:0] MemController_34_io_rd_data_bits; // @[pearray.scala 200:15]
  wire  MemController_34_io_wr_data_valid; // @[pearray.scala 200:15]
  wire [7:0] MemController_34_io_wr_data_bits; // @[pearray.scala 200:15]
  wire  MemController_35_clock; // @[pearray.scala 200:15]
  wire  MemController_35_reset; // @[pearray.scala 200:15]
  wire  MemController_35_io_rd_valid; // @[pearray.scala 200:15]
  wire  MemController_35_io_wr_valid; // @[pearray.scala 200:15]
  wire  MemController_35_io_rd_data_valid; // @[pearray.scala 200:15]
  wire [7:0] MemController_35_io_rd_data_bits; // @[pearray.scala 200:15]
  wire  MemController_35_io_wr_data_valid; // @[pearray.scala 200:15]
  wire [7:0] MemController_35_io_wr_data_bits; // @[pearray.scala 200:15]
  wire  MemController_36_clock; // @[pearray.scala 200:15]
  wire  MemController_36_reset; // @[pearray.scala 200:15]
  wire  MemController_36_io_rd_valid; // @[pearray.scala 200:15]
  wire  MemController_36_io_wr_valid; // @[pearray.scala 200:15]
  wire  MemController_36_io_rd_data_valid; // @[pearray.scala 200:15]
  wire [7:0] MemController_36_io_rd_data_bits; // @[pearray.scala 200:15]
  wire  MemController_36_io_wr_data_valid; // @[pearray.scala 200:15]
  wire [7:0] MemController_36_io_wr_data_bits; // @[pearray.scala 200:15]
  wire  MemController_37_clock; // @[pearray.scala 200:15]
  wire  MemController_37_reset; // @[pearray.scala 200:15]
  wire  MemController_37_io_rd_valid; // @[pearray.scala 200:15]
  wire  MemController_37_io_wr_valid; // @[pearray.scala 200:15]
  wire  MemController_37_io_rd_data_valid; // @[pearray.scala 200:15]
  wire [7:0] MemController_37_io_rd_data_bits; // @[pearray.scala 200:15]
  wire  MemController_37_io_wr_data_valid; // @[pearray.scala 200:15]
  wire [7:0] MemController_37_io_wr_data_bits; // @[pearray.scala 200:15]
  wire  MemController_38_clock; // @[pearray.scala 200:15]
  wire  MemController_38_reset; // @[pearray.scala 200:15]
  wire  MemController_38_io_rd_valid; // @[pearray.scala 200:15]
  wire  MemController_38_io_wr_valid; // @[pearray.scala 200:15]
  wire  MemController_38_io_rd_data_valid; // @[pearray.scala 200:15]
  wire [7:0] MemController_38_io_rd_data_bits; // @[pearray.scala 200:15]
  wire  MemController_38_io_wr_data_valid; // @[pearray.scala 200:15]
  wire [7:0] MemController_38_io_wr_data_bits; // @[pearray.scala 200:15]
  wire  MemController_39_clock; // @[pearray.scala 200:15]
  wire  MemController_39_reset; // @[pearray.scala 200:15]
  wire  MemController_39_io_rd_valid; // @[pearray.scala 200:15]
  wire  MemController_39_io_wr_valid; // @[pearray.scala 200:15]
  wire  MemController_39_io_rd_data_valid; // @[pearray.scala 200:15]
  wire [7:0] MemController_39_io_rd_data_bits; // @[pearray.scala 200:15]
  wire  MemController_39_io_wr_data_valid; // @[pearray.scala 200:15]
  wire [7:0] MemController_39_io_wr_data_bits; // @[pearray.scala 200:15]
  wire  _T_1 = ~reset; // @[pearray.scala 64:9]
  wire  _T_7 = MultiDimTime_io_index_1 == 18'h0; // @[pearray.scala 180:73]
  wire  _T_8 = MultiDimTime_io_index_0 == 18'h0; // @[pearray.scala 180:121]
  wire  _T_9 = _T_7 & _T_8; // @[pearray.scala 180:99]
  reg  _T_16_0; // @[pearray.scala 51:27]
  reg [31:0] _RAND_0;
  reg  _T_16_1; // @[pearray.scala 51:27]
  reg [31:0] _RAND_1;
  reg  _T_16_2; // @[pearray.scala 51:27]
  reg [31:0] _RAND_2;
  reg  _T_16_3; // @[pearray.scala 51:27]
  reg [31:0] _RAND_3;
  wire  _T_19 = MultiDimTime_io_index_1 == 18'h1; // @[pearray.scala 180:73]
  wire  _T_21 = _T_19 & _T_8; // @[pearray.scala 180:99]
  reg  _T_28_0; // @[pearray.scala 51:27]
  reg [31:0] _RAND_4;
  reg  _T_28_1; // @[pearray.scala 51:27]
  reg [31:0] _RAND_5;
  reg  _T_28_2; // @[pearray.scala 51:27]
  reg [31:0] _RAND_6;
  reg  _T_28_3; // @[pearray.scala 51:27]
  reg [31:0] _RAND_7;
  wire  _T_31 = MultiDimTime_io_index_1 == 18'h2; // @[pearray.scala 180:73]
  wire  _T_33 = _T_31 & _T_8; // @[pearray.scala 180:99]
  reg  _T_40_0; // @[pearray.scala 51:27]
  reg [31:0] _RAND_8;
  reg  _T_40_1; // @[pearray.scala 51:27]
  reg [31:0] _RAND_9;
  reg  _T_40_2; // @[pearray.scala 51:27]
  reg [31:0] _RAND_10;
  reg  _T_40_3; // @[pearray.scala 51:27]
  reg [31:0] _RAND_11;
  wire  _T_43 = MultiDimTime_io_index_1 == 18'h3; // @[pearray.scala 180:73]
  wire  _T_45 = _T_43 & _T_8; // @[pearray.scala 180:99]
  reg  _T_52_0; // @[pearray.scala 51:27]
  reg [31:0] _RAND_12;
  reg  _T_52_1; // @[pearray.scala 51:27]
  reg [31:0] _RAND_13;
  reg  _T_52_2; // @[pearray.scala 51:27]
  reg [31:0] _RAND_14;
  reg  _T_52_3; // @[pearray.scala 51:27]
  reg [31:0] _RAND_15;
  wire  _T_55 = MultiDimTime_io_index_1 == 18'h4; // @[pearray.scala 180:73]
  wire  _T_57 = _T_55 & _T_8; // @[pearray.scala 180:99]
  reg  _T_64_0; // @[pearray.scala 51:27]
  reg [31:0] _RAND_16;
  reg  _T_64_1; // @[pearray.scala 51:27]
  reg [31:0] _RAND_17;
  reg  _T_64_2; // @[pearray.scala 51:27]
  reg [31:0] _RAND_18;
  reg  _T_64_3; // @[pearray.scala 51:27]
  reg [31:0] _RAND_19;
  wire  _T_67 = MultiDimTime_io_index_1 == 18'h5; // @[pearray.scala 180:73]
  wire  _T_69 = _T_67 & _T_8; // @[pearray.scala 180:99]
  reg  _T_76_0; // @[pearray.scala 51:27]
  reg [31:0] _RAND_20;
  reg  _T_76_1; // @[pearray.scala 51:27]
  reg [31:0] _RAND_21;
  reg  _T_76_2; // @[pearray.scala 51:27]
  reg [31:0] _RAND_22;
  reg  _T_76_3; // @[pearray.scala 51:27]
  reg [31:0] _RAND_23;
  wire  _T_79 = MultiDimTime_io_index_1 == 18'h6; // @[pearray.scala 180:73]
  wire  _T_81 = _T_79 & _T_8; // @[pearray.scala 180:99]
  reg  _T_88_0; // @[pearray.scala 51:27]
  reg [31:0] _RAND_24;
  reg  _T_88_1; // @[pearray.scala 51:27]
  reg [31:0] _RAND_25;
  reg  _T_88_2; // @[pearray.scala 51:27]
  reg [31:0] _RAND_26;
  reg  _T_88_3; // @[pearray.scala 51:27]
  reg [31:0] _RAND_27;
  wire  _T_91 = MultiDimTime_io_index_1 == 18'h7; // @[pearray.scala 180:73]
  wire  _T_93 = _T_91 & _T_8; // @[pearray.scala 180:99]
  reg  _T_100_0; // @[pearray.scala 51:27]
  reg [31:0] _RAND_28;
  reg  _T_100_1; // @[pearray.scala 51:27]
  reg [31:0] _RAND_29;
  reg  _T_100_2; // @[pearray.scala 51:27]
  reg [31:0] _RAND_30;
  reg  _T_100_3; // @[pearray.scala 51:27]
  reg [31:0] _RAND_31;
  reg  _T_114_0; // @[pearray.scala 51:27]
  reg [31:0] _RAND_32;
  reg  _T_114_1; // @[pearray.scala 51:27]
  reg [31:0] _RAND_33;
  reg  _T_114_2; // @[pearray.scala 51:27]
  reg [31:0] _RAND_34;
  reg  _T_114_3; // @[pearray.scala 51:27]
  reg [31:0] _RAND_35;
  reg  _T_126_0; // @[pearray.scala 51:27]
  reg [31:0] _RAND_36;
  reg  _T_126_1; // @[pearray.scala 51:27]
  reg [31:0] _RAND_37;
  reg  _T_126_2; // @[pearray.scala 51:27]
  reg [31:0] _RAND_38;
  reg  _T_126_3; // @[pearray.scala 51:27]
  reg [31:0] _RAND_39;
  reg  _T_138_0; // @[pearray.scala 51:27]
  reg [31:0] _RAND_40;
  reg  _T_138_1; // @[pearray.scala 51:27]
  reg [31:0] _RAND_41;
  reg  _T_138_2; // @[pearray.scala 51:27]
  reg [31:0] _RAND_42;
  reg  _T_138_3; // @[pearray.scala 51:27]
  reg [31:0] _RAND_43;
  reg  _T_150_0; // @[pearray.scala 51:27]
  reg [31:0] _RAND_44;
  reg  _T_150_1; // @[pearray.scala 51:27]
  reg [31:0] _RAND_45;
  reg  _T_150_2; // @[pearray.scala 51:27]
  reg [31:0] _RAND_46;
  reg  _T_150_3; // @[pearray.scala 51:27]
  reg [31:0] _RAND_47;
  reg  _T_162_0; // @[pearray.scala 51:27]
  reg [31:0] _RAND_48;
  reg  _T_162_1; // @[pearray.scala 51:27]
  reg [31:0] _RAND_49;
  reg  _T_162_2; // @[pearray.scala 51:27]
  reg [31:0] _RAND_50;
  reg  _T_162_3; // @[pearray.scala 51:27]
  reg [31:0] _RAND_51;
  reg  _T_174_0; // @[pearray.scala 51:27]
  reg [31:0] _RAND_52;
  reg  _T_174_1; // @[pearray.scala 51:27]
  reg [31:0] _RAND_53;
  reg  _T_174_2; // @[pearray.scala 51:27]
  reg [31:0] _RAND_54;
  reg  _T_174_3; // @[pearray.scala 51:27]
  reg [31:0] _RAND_55;
  reg  _T_186_0; // @[pearray.scala 51:27]
  reg [31:0] _RAND_56;
  reg  _T_186_1; // @[pearray.scala 51:27]
  reg [31:0] _RAND_57;
  reg  _T_186_2; // @[pearray.scala 51:27]
  reg [31:0] _RAND_58;
  reg  _T_186_3; // @[pearray.scala 51:27]
  reg [31:0] _RAND_59;
  wire  _T_189 = MultiDimTime_io_index_1 == 18'h8; // @[pearray.scala 180:73]
  wire  _T_191 = _T_189 & _T_8; // @[pearray.scala 180:99]
  reg  _T_198_0; // @[pearray.scala 51:27]
  reg [31:0] _RAND_60;
  reg  _T_198_1; // @[pearray.scala 51:27]
  reg [31:0] _RAND_61;
  reg  _T_198_2; // @[pearray.scala 51:27]
  reg [31:0] _RAND_62;
  reg  _T_198_3; // @[pearray.scala 51:27]
  reg [31:0] _RAND_63;
  reg  _T_212_0; // @[pearray.scala 51:27]
  reg [31:0] _RAND_64;
  reg  _T_212_1; // @[pearray.scala 51:27]
  reg [31:0] _RAND_65;
  reg  _T_212_2; // @[pearray.scala 51:27]
  reg [31:0] _RAND_66;
  reg  _T_212_3; // @[pearray.scala 51:27]
  reg [31:0] _RAND_67;
  reg  _T_224_0; // @[pearray.scala 51:27]
  reg [31:0] _RAND_68;
  reg  _T_224_1; // @[pearray.scala 51:27]
  reg [31:0] _RAND_69;
  reg  _T_224_2; // @[pearray.scala 51:27]
  reg [31:0] _RAND_70;
  reg  _T_224_3; // @[pearray.scala 51:27]
  reg [31:0] _RAND_71;
  reg  _T_236_0; // @[pearray.scala 51:27]
  reg [31:0] _RAND_72;
  reg  _T_236_1; // @[pearray.scala 51:27]
  reg [31:0] _RAND_73;
  reg  _T_236_2; // @[pearray.scala 51:27]
  reg [31:0] _RAND_74;
  reg  _T_236_3; // @[pearray.scala 51:27]
  reg [31:0] _RAND_75;
  reg  _T_248_0; // @[pearray.scala 51:27]
  reg [31:0] _RAND_76;
  reg  _T_248_1; // @[pearray.scala 51:27]
  reg [31:0] _RAND_77;
  reg  _T_248_2; // @[pearray.scala 51:27]
  reg [31:0] _RAND_78;
  reg  _T_248_3; // @[pearray.scala 51:27]
  reg [31:0] _RAND_79;
  reg  _T_260_0; // @[pearray.scala 51:27]
  reg [31:0] _RAND_80;
  reg  _T_260_1; // @[pearray.scala 51:27]
  reg [31:0] _RAND_81;
  reg  _T_260_2; // @[pearray.scala 51:27]
  reg [31:0] _RAND_82;
  reg  _T_260_3; // @[pearray.scala 51:27]
  reg [31:0] _RAND_83;
  reg  _T_272_0; // @[pearray.scala 51:27]
  reg [31:0] _RAND_84;
  reg  _T_272_1; // @[pearray.scala 51:27]
  reg [31:0] _RAND_85;
  reg  _T_272_2; // @[pearray.scala 51:27]
  reg [31:0] _RAND_86;
  reg  _T_272_3; // @[pearray.scala 51:27]
  reg [31:0] _RAND_87;
  reg  _T_284_0; // @[pearray.scala 51:27]
  reg [31:0] _RAND_88;
  reg  _T_284_1; // @[pearray.scala 51:27]
  reg [31:0] _RAND_89;
  reg  _T_284_2; // @[pearray.scala 51:27]
  reg [31:0] _RAND_90;
  reg  _T_284_3; // @[pearray.scala 51:27]
  reg [31:0] _RAND_91;
  wire  _T_287 = MultiDimTime_io_index_1 == 18'h9; // @[pearray.scala 180:73]
  wire  _T_289 = _T_287 & _T_8; // @[pearray.scala 180:99]
  reg  _T_296_0; // @[pearray.scala 51:27]
  reg [31:0] _RAND_92;
  reg  _T_296_1; // @[pearray.scala 51:27]
  reg [31:0] _RAND_93;
  reg  _T_296_2; // @[pearray.scala 51:27]
  reg [31:0] _RAND_94;
  reg  _T_296_3; // @[pearray.scala 51:27]
  reg [31:0] _RAND_95;
  reg  _T_310_0; // @[pearray.scala 51:27]
  reg [31:0] _RAND_96;
  reg  _T_310_1; // @[pearray.scala 51:27]
  reg [31:0] _RAND_97;
  reg  _T_310_2; // @[pearray.scala 51:27]
  reg [31:0] _RAND_98;
  reg  _T_310_3; // @[pearray.scala 51:27]
  reg [31:0] _RAND_99;
  reg  _T_322_0; // @[pearray.scala 51:27]
  reg [31:0] _RAND_100;
  reg  _T_322_1; // @[pearray.scala 51:27]
  reg [31:0] _RAND_101;
  reg  _T_322_2; // @[pearray.scala 51:27]
  reg [31:0] _RAND_102;
  reg  _T_322_3; // @[pearray.scala 51:27]
  reg [31:0] _RAND_103;
  reg  _T_334_0; // @[pearray.scala 51:27]
  reg [31:0] _RAND_104;
  reg  _T_334_1; // @[pearray.scala 51:27]
  reg [31:0] _RAND_105;
  reg  _T_334_2; // @[pearray.scala 51:27]
  reg [31:0] _RAND_106;
  reg  _T_334_3; // @[pearray.scala 51:27]
  reg [31:0] _RAND_107;
  reg  _T_346_0; // @[pearray.scala 51:27]
  reg [31:0] _RAND_108;
  reg  _T_346_1; // @[pearray.scala 51:27]
  reg [31:0] _RAND_109;
  reg  _T_346_2; // @[pearray.scala 51:27]
  reg [31:0] _RAND_110;
  reg  _T_346_3; // @[pearray.scala 51:27]
  reg [31:0] _RAND_111;
  reg  _T_358_0; // @[pearray.scala 51:27]
  reg [31:0] _RAND_112;
  reg  _T_358_1; // @[pearray.scala 51:27]
  reg [31:0] _RAND_113;
  reg  _T_358_2; // @[pearray.scala 51:27]
  reg [31:0] _RAND_114;
  reg  _T_358_3; // @[pearray.scala 51:27]
  reg [31:0] _RAND_115;
  reg  _T_370_0; // @[pearray.scala 51:27]
  reg [31:0] _RAND_116;
  reg  _T_370_1; // @[pearray.scala 51:27]
  reg [31:0] _RAND_117;
  reg  _T_370_2; // @[pearray.scala 51:27]
  reg [31:0] _RAND_118;
  reg  _T_370_3; // @[pearray.scala 51:27]
  reg [31:0] _RAND_119;
  reg  _T_382_0; // @[pearray.scala 51:27]
  reg [31:0] _RAND_120;
  reg  _T_382_1; // @[pearray.scala 51:27]
  reg [31:0] _RAND_121;
  reg  _T_382_2; // @[pearray.scala 51:27]
  reg [31:0] _RAND_122;
  reg  _T_382_3; // @[pearray.scala 51:27]
  reg [31:0] _RAND_123;
  wire  _T_385 = MultiDimTime_io_index_1 == 18'ha; // @[pearray.scala 180:73]
  wire  _T_387 = _T_385 & _T_8; // @[pearray.scala 180:99]
  reg  _T_394_0; // @[pearray.scala 51:27]
  reg [31:0] _RAND_124;
  reg  _T_394_1; // @[pearray.scala 51:27]
  reg [31:0] _RAND_125;
  reg  _T_394_2; // @[pearray.scala 51:27]
  reg [31:0] _RAND_126;
  reg  _T_394_3; // @[pearray.scala 51:27]
  reg [31:0] _RAND_127;
  reg  _T_408_0; // @[pearray.scala 51:27]
  reg [31:0] _RAND_128;
  reg  _T_408_1; // @[pearray.scala 51:27]
  reg [31:0] _RAND_129;
  reg  _T_408_2; // @[pearray.scala 51:27]
  reg [31:0] _RAND_130;
  reg  _T_408_3; // @[pearray.scala 51:27]
  reg [31:0] _RAND_131;
  reg  _T_420_0; // @[pearray.scala 51:27]
  reg [31:0] _RAND_132;
  reg  _T_420_1; // @[pearray.scala 51:27]
  reg [31:0] _RAND_133;
  reg  _T_420_2; // @[pearray.scala 51:27]
  reg [31:0] _RAND_134;
  reg  _T_420_3; // @[pearray.scala 51:27]
  reg [31:0] _RAND_135;
  reg  _T_432_0; // @[pearray.scala 51:27]
  reg [31:0] _RAND_136;
  reg  _T_432_1; // @[pearray.scala 51:27]
  reg [31:0] _RAND_137;
  reg  _T_432_2; // @[pearray.scala 51:27]
  reg [31:0] _RAND_138;
  reg  _T_432_3; // @[pearray.scala 51:27]
  reg [31:0] _RAND_139;
  reg  _T_444_0; // @[pearray.scala 51:27]
  reg [31:0] _RAND_140;
  reg  _T_444_1; // @[pearray.scala 51:27]
  reg [31:0] _RAND_141;
  reg  _T_444_2; // @[pearray.scala 51:27]
  reg [31:0] _RAND_142;
  reg  _T_444_3; // @[pearray.scala 51:27]
  reg [31:0] _RAND_143;
  reg  _T_456_0; // @[pearray.scala 51:27]
  reg [31:0] _RAND_144;
  reg  _T_456_1; // @[pearray.scala 51:27]
  reg [31:0] _RAND_145;
  reg  _T_456_2; // @[pearray.scala 51:27]
  reg [31:0] _RAND_146;
  reg  _T_456_3; // @[pearray.scala 51:27]
  reg [31:0] _RAND_147;
  reg  _T_468_0; // @[pearray.scala 51:27]
  reg [31:0] _RAND_148;
  reg  _T_468_1; // @[pearray.scala 51:27]
  reg [31:0] _RAND_149;
  reg  _T_468_2; // @[pearray.scala 51:27]
  reg [31:0] _RAND_150;
  reg  _T_468_3; // @[pearray.scala 51:27]
  reg [31:0] _RAND_151;
  reg  _T_480_0; // @[pearray.scala 51:27]
  reg [31:0] _RAND_152;
  reg  _T_480_1; // @[pearray.scala 51:27]
  reg [31:0] _RAND_153;
  reg  _T_480_2; // @[pearray.scala 51:27]
  reg [31:0] _RAND_154;
  reg  _T_480_3; // @[pearray.scala 51:27]
  reg [31:0] _RAND_155;
  wire  _T_483 = MultiDimTime_io_index_1 == 18'hb; // @[pearray.scala 180:73]
  wire  _T_485 = _T_483 & _T_8; // @[pearray.scala 180:99]
  reg  _T_492_0; // @[pearray.scala 51:27]
  reg [31:0] _RAND_156;
  reg  _T_492_1; // @[pearray.scala 51:27]
  reg [31:0] _RAND_157;
  reg  _T_492_2; // @[pearray.scala 51:27]
  reg [31:0] _RAND_158;
  reg  _T_492_3; // @[pearray.scala 51:27]
  reg [31:0] _RAND_159;
  reg  _T_506_0; // @[pearray.scala 51:27]
  reg [31:0] _RAND_160;
  reg  _T_506_1; // @[pearray.scala 51:27]
  reg [31:0] _RAND_161;
  reg  _T_506_2; // @[pearray.scala 51:27]
  reg [31:0] _RAND_162;
  reg  _T_506_3; // @[pearray.scala 51:27]
  reg [31:0] _RAND_163;
  reg  _T_518_0; // @[pearray.scala 51:27]
  reg [31:0] _RAND_164;
  reg  _T_518_1; // @[pearray.scala 51:27]
  reg [31:0] _RAND_165;
  reg  _T_518_2; // @[pearray.scala 51:27]
  reg [31:0] _RAND_166;
  reg  _T_518_3; // @[pearray.scala 51:27]
  reg [31:0] _RAND_167;
  reg  _T_530_0; // @[pearray.scala 51:27]
  reg [31:0] _RAND_168;
  reg  _T_530_1; // @[pearray.scala 51:27]
  reg [31:0] _RAND_169;
  reg  _T_530_2; // @[pearray.scala 51:27]
  reg [31:0] _RAND_170;
  reg  _T_530_3; // @[pearray.scala 51:27]
  reg [31:0] _RAND_171;
  reg  _T_542_0; // @[pearray.scala 51:27]
  reg [31:0] _RAND_172;
  reg  _T_542_1; // @[pearray.scala 51:27]
  reg [31:0] _RAND_173;
  reg  _T_542_2; // @[pearray.scala 51:27]
  reg [31:0] _RAND_174;
  reg  _T_542_3; // @[pearray.scala 51:27]
  reg [31:0] _RAND_175;
  reg  _T_554_0; // @[pearray.scala 51:27]
  reg [31:0] _RAND_176;
  reg  _T_554_1; // @[pearray.scala 51:27]
  reg [31:0] _RAND_177;
  reg  _T_554_2; // @[pearray.scala 51:27]
  reg [31:0] _RAND_178;
  reg  _T_554_3; // @[pearray.scala 51:27]
  reg [31:0] _RAND_179;
  reg  _T_566_0; // @[pearray.scala 51:27]
  reg [31:0] _RAND_180;
  reg  _T_566_1; // @[pearray.scala 51:27]
  reg [31:0] _RAND_181;
  reg  _T_566_2; // @[pearray.scala 51:27]
  reg [31:0] _RAND_182;
  reg  _T_566_3; // @[pearray.scala 51:27]
  reg [31:0] _RAND_183;
  reg  _T_578_0; // @[pearray.scala 51:27]
  reg [31:0] _RAND_184;
  reg  _T_578_1; // @[pearray.scala 51:27]
  reg [31:0] _RAND_185;
  reg  _T_578_2; // @[pearray.scala 51:27]
  reg [31:0] _RAND_186;
  reg  _T_578_3; // @[pearray.scala 51:27]
  reg [31:0] _RAND_187;
  wire  _T_581 = MultiDimTime_io_index_1 == 18'hc; // @[pearray.scala 180:73]
  wire  _T_583 = _T_581 & _T_8; // @[pearray.scala 180:99]
  reg  _T_590_0; // @[pearray.scala 51:27]
  reg [31:0] _RAND_188;
  reg  _T_590_1; // @[pearray.scala 51:27]
  reg [31:0] _RAND_189;
  reg  _T_590_2; // @[pearray.scala 51:27]
  reg [31:0] _RAND_190;
  reg  _T_590_3; // @[pearray.scala 51:27]
  reg [31:0] _RAND_191;
  reg  _T_604_0; // @[pearray.scala 51:27]
  reg [31:0] _RAND_192;
  reg  _T_604_1; // @[pearray.scala 51:27]
  reg [31:0] _RAND_193;
  reg  _T_604_2; // @[pearray.scala 51:27]
  reg [31:0] _RAND_194;
  reg  _T_604_3; // @[pearray.scala 51:27]
  reg [31:0] _RAND_195;
  reg  _T_616_0; // @[pearray.scala 51:27]
  reg [31:0] _RAND_196;
  reg  _T_616_1; // @[pearray.scala 51:27]
  reg [31:0] _RAND_197;
  reg  _T_616_2; // @[pearray.scala 51:27]
  reg [31:0] _RAND_198;
  reg  _T_616_3; // @[pearray.scala 51:27]
  reg [31:0] _RAND_199;
  reg  _T_628_0; // @[pearray.scala 51:27]
  reg [31:0] _RAND_200;
  reg  _T_628_1; // @[pearray.scala 51:27]
  reg [31:0] _RAND_201;
  reg  _T_628_2; // @[pearray.scala 51:27]
  reg [31:0] _RAND_202;
  reg  _T_628_3; // @[pearray.scala 51:27]
  reg [31:0] _RAND_203;
  reg  _T_640_0; // @[pearray.scala 51:27]
  reg [31:0] _RAND_204;
  reg  _T_640_1; // @[pearray.scala 51:27]
  reg [31:0] _RAND_205;
  reg  _T_640_2; // @[pearray.scala 51:27]
  reg [31:0] _RAND_206;
  reg  _T_640_3; // @[pearray.scala 51:27]
  reg [31:0] _RAND_207;
  reg  _T_652_0; // @[pearray.scala 51:27]
  reg [31:0] _RAND_208;
  reg  _T_652_1; // @[pearray.scala 51:27]
  reg [31:0] _RAND_209;
  reg  _T_652_2; // @[pearray.scala 51:27]
  reg [31:0] _RAND_210;
  reg  _T_652_3; // @[pearray.scala 51:27]
  reg [31:0] _RAND_211;
  reg  _T_664_0; // @[pearray.scala 51:27]
  reg [31:0] _RAND_212;
  reg  _T_664_1; // @[pearray.scala 51:27]
  reg [31:0] _RAND_213;
  reg  _T_664_2; // @[pearray.scala 51:27]
  reg [31:0] _RAND_214;
  reg  _T_664_3; // @[pearray.scala 51:27]
  reg [31:0] _RAND_215;
  reg  _T_676_0; // @[pearray.scala 51:27]
  reg [31:0] _RAND_216;
  reg  _T_676_1; // @[pearray.scala 51:27]
  reg [31:0] _RAND_217;
  reg  _T_676_2; // @[pearray.scala 51:27]
  reg [31:0] _RAND_218;
  reg  _T_676_3; // @[pearray.scala 51:27]
  reg [31:0] _RAND_219;
  wire  _T_679 = MultiDimTime_io_index_1 == 18'hd; // @[pearray.scala 180:73]
  wire  _T_681 = _T_679 & _T_8; // @[pearray.scala 180:99]
  reg  _T_688_0; // @[pearray.scala 51:27]
  reg [31:0] _RAND_220;
  reg  _T_688_1; // @[pearray.scala 51:27]
  reg [31:0] _RAND_221;
  reg  _T_688_2; // @[pearray.scala 51:27]
  reg [31:0] _RAND_222;
  reg  _T_688_3; // @[pearray.scala 51:27]
  reg [31:0] _RAND_223;
  reg  _T_702_0; // @[pearray.scala 51:27]
  reg [31:0] _RAND_224;
  reg  _T_702_1; // @[pearray.scala 51:27]
  reg [31:0] _RAND_225;
  reg  _T_702_2; // @[pearray.scala 51:27]
  reg [31:0] _RAND_226;
  reg  _T_702_3; // @[pearray.scala 51:27]
  reg [31:0] _RAND_227;
  reg  _T_714_0; // @[pearray.scala 51:27]
  reg [31:0] _RAND_228;
  reg  _T_714_1; // @[pearray.scala 51:27]
  reg [31:0] _RAND_229;
  reg  _T_714_2; // @[pearray.scala 51:27]
  reg [31:0] _RAND_230;
  reg  _T_714_3; // @[pearray.scala 51:27]
  reg [31:0] _RAND_231;
  reg  _T_726_0; // @[pearray.scala 51:27]
  reg [31:0] _RAND_232;
  reg  _T_726_1; // @[pearray.scala 51:27]
  reg [31:0] _RAND_233;
  reg  _T_726_2; // @[pearray.scala 51:27]
  reg [31:0] _RAND_234;
  reg  _T_726_3; // @[pearray.scala 51:27]
  reg [31:0] _RAND_235;
  reg  _T_738_0; // @[pearray.scala 51:27]
  reg [31:0] _RAND_236;
  reg  _T_738_1; // @[pearray.scala 51:27]
  reg [31:0] _RAND_237;
  reg  _T_738_2; // @[pearray.scala 51:27]
  reg [31:0] _RAND_238;
  reg  _T_738_3; // @[pearray.scala 51:27]
  reg [31:0] _RAND_239;
  reg  _T_750_0; // @[pearray.scala 51:27]
  reg [31:0] _RAND_240;
  reg  _T_750_1; // @[pearray.scala 51:27]
  reg [31:0] _RAND_241;
  reg  _T_750_2; // @[pearray.scala 51:27]
  reg [31:0] _RAND_242;
  reg  _T_750_3; // @[pearray.scala 51:27]
  reg [31:0] _RAND_243;
  reg  _T_762_0; // @[pearray.scala 51:27]
  reg [31:0] _RAND_244;
  reg  _T_762_1; // @[pearray.scala 51:27]
  reg [31:0] _RAND_245;
  reg  _T_762_2; // @[pearray.scala 51:27]
  reg [31:0] _RAND_246;
  reg  _T_762_3; // @[pearray.scala 51:27]
  reg [31:0] _RAND_247;
  reg  _T_774_0; // @[pearray.scala 51:27]
  reg [31:0] _RAND_248;
  reg  _T_774_1; // @[pearray.scala 51:27]
  reg [31:0] _RAND_249;
  reg  _T_774_2; // @[pearray.scala 51:27]
  reg [31:0] _RAND_250;
  reg  _T_774_3; // @[pearray.scala 51:27]
  reg [31:0] _RAND_251;
  wire  _T_777 = MultiDimTime_io_index_1 == 18'he; // @[pearray.scala 180:73]
  wire  _T_779 = _T_777 & _T_8; // @[pearray.scala 180:99]
  reg  _T_786_0; // @[pearray.scala 51:27]
  reg [31:0] _RAND_252;
  reg  _T_786_1; // @[pearray.scala 51:27]
  reg [31:0] _RAND_253;
  reg  _T_786_2; // @[pearray.scala 51:27]
  reg [31:0] _RAND_254;
  reg  _T_786_3; // @[pearray.scala 51:27]
  reg [31:0] _RAND_255;
  reg  _T_800_0; // @[pearray.scala 51:27]
  reg [31:0] _RAND_256;
  reg  _T_800_1; // @[pearray.scala 51:27]
  reg [31:0] _RAND_257;
  reg  _T_800_2; // @[pearray.scala 51:27]
  reg [31:0] _RAND_258;
  reg  _T_800_3; // @[pearray.scala 51:27]
  reg [31:0] _RAND_259;
  reg  _T_812_0; // @[pearray.scala 51:27]
  reg [31:0] _RAND_260;
  reg  _T_812_1; // @[pearray.scala 51:27]
  reg [31:0] _RAND_261;
  reg  _T_812_2; // @[pearray.scala 51:27]
  reg [31:0] _RAND_262;
  reg  _T_812_3; // @[pearray.scala 51:27]
  reg [31:0] _RAND_263;
  reg  _T_824_0; // @[pearray.scala 51:27]
  reg [31:0] _RAND_264;
  reg  _T_824_1; // @[pearray.scala 51:27]
  reg [31:0] _RAND_265;
  reg  _T_824_2; // @[pearray.scala 51:27]
  reg [31:0] _RAND_266;
  reg  _T_824_3; // @[pearray.scala 51:27]
  reg [31:0] _RAND_267;
  reg  _T_836_0; // @[pearray.scala 51:27]
  reg [31:0] _RAND_268;
  reg  _T_836_1; // @[pearray.scala 51:27]
  reg [31:0] _RAND_269;
  reg  _T_836_2; // @[pearray.scala 51:27]
  reg [31:0] _RAND_270;
  reg  _T_836_3; // @[pearray.scala 51:27]
  reg [31:0] _RAND_271;
  reg  _T_848_0; // @[pearray.scala 51:27]
  reg [31:0] _RAND_272;
  reg  _T_848_1; // @[pearray.scala 51:27]
  reg [31:0] _RAND_273;
  reg  _T_848_2; // @[pearray.scala 51:27]
  reg [31:0] _RAND_274;
  reg  _T_848_3; // @[pearray.scala 51:27]
  reg [31:0] _RAND_275;
  reg  _T_860_0; // @[pearray.scala 51:27]
  reg [31:0] _RAND_276;
  reg  _T_860_1; // @[pearray.scala 51:27]
  reg [31:0] _RAND_277;
  reg  _T_860_2; // @[pearray.scala 51:27]
  reg [31:0] _RAND_278;
  reg  _T_860_3; // @[pearray.scala 51:27]
  reg [31:0] _RAND_279;
  reg  _T_872_0; // @[pearray.scala 51:27]
  reg [31:0] _RAND_280;
  reg  _T_872_1; // @[pearray.scala 51:27]
  reg [31:0] _RAND_281;
  reg  _T_872_2; // @[pearray.scala 51:27]
  reg [31:0] _RAND_282;
  reg  _T_872_3; // @[pearray.scala 51:27]
  reg [31:0] _RAND_283;
  wire  _T_875 = MultiDimTime_io_index_1 == 18'hf; // @[pearray.scala 180:73]
  wire  _T_877 = _T_875 & _T_8; // @[pearray.scala 180:99]
  reg  _T_884_0; // @[pearray.scala 51:27]
  reg [31:0] _RAND_284;
  reg  _T_884_1; // @[pearray.scala 51:27]
  reg [31:0] _RAND_285;
  reg  _T_884_2; // @[pearray.scala 51:27]
  reg [31:0] _RAND_286;
  reg  _T_884_3; // @[pearray.scala 51:27]
  reg [31:0] _RAND_287;
  reg  _T_898_0; // @[pearray.scala 51:27]
  reg [31:0] _RAND_288;
  reg  _T_898_1; // @[pearray.scala 51:27]
  reg [31:0] _RAND_289;
  reg  _T_898_2; // @[pearray.scala 51:27]
  reg [31:0] _RAND_290;
  reg  _T_898_3; // @[pearray.scala 51:27]
  reg [31:0] _RAND_291;
  reg  _T_910_0; // @[pearray.scala 51:27]
  reg [31:0] _RAND_292;
  reg  _T_910_1; // @[pearray.scala 51:27]
  reg [31:0] _RAND_293;
  reg  _T_910_2; // @[pearray.scala 51:27]
  reg [31:0] _RAND_294;
  reg  _T_910_3; // @[pearray.scala 51:27]
  reg [31:0] _RAND_295;
  reg  _T_922_0; // @[pearray.scala 51:27]
  reg [31:0] _RAND_296;
  reg  _T_922_1; // @[pearray.scala 51:27]
  reg [31:0] _RAND_297;
  reg  _T_922_2; // @[pearray.scala 51:27]
  reg [31:0] _RAND_298;
  reg  _T_922_3; // @[pearray.scala 51:27]
  reg [31:0] _RAND_299;
  reg  _T_934_0; // @[pearray.scala 51:27]
  reg [31:0] _RAND_300;
  reg  _T_934_1; // @[pearray.scala 51:27]
  reg [31:0] _RAND_301;
  reg  _T_934_2; // @[pearray.scala 51:27]
  reg [31:0] _RAND_302;
  reg  _T_934_3; // @[pearray.scala 51:27]
  reg [31:0] _RAND_303;
  reg  _T_946_0; // @[pearray.scala 51:27]
  reg [31:0] _RAND_304;
  reg  _T_946_1; // @[pearray.scala 51:27]
  reg [31:0] _RAND_305;
  reg  _T_946_2; // @[pearray.scala 51:27]
  reg [31:0] _RAND_306;
  reg  _T_946_3; // @[pearray.scala 51:27]
  reg [31:0] _RAND_307;
  reg  _T_958_0; // @[pearray.scala 51:27]
  reg [31:0] _RAND_308;
  reg  _T_958_1; // @[pearray.scala 51:27]
  reg [31:0] _RAND_309;
  reg  _T_958_2; // @[pearray.scala 51:27]
  reg [31:0] _RAND_310;
  reg  _T_958_3; // @[pearray.scala 51:27]
  reg [31:0] _RAND_311;
  reg  _T_970_0; // @[pearray.scala 51:27]
  reg [31:0] _RAND_312;
  reg  _T_970_1; // @[pearray.scala 51:27]
  reg [31:0] _RAND_313;
  reg  _T_970_2; // @[pearray.scala 51:27]
  reg [31:0] _RAND_314;
  reg  _T_970_3; // @[pearray.scala 51:27]
  reg [31:0] _RAND_315;
  wire  _T_973 = MultiDimTime_io_index_1 == 18'h10; // @[pearray.scala 180:73]
  wire  _T_975 = _T_973 & _T_8; // @[pearray.scala 180:99]
  reg  _T_982_0; // @[pearray.scala 51:27]
  reg [31:0] _RAND_316;
  reg  _T_982_1; // @[pearray.scala 51:27]
  reg [31:0] _RAND_317;
  reg  _T_982_2; // @[pearray.scala 51:27]
  reg [31:0] _RAND_318;
  reg  _T_982_3; // @[pearray.scala 51:27]
  reg [31:0] _RAND_319;
  reg  _T_996_0; // @[pearray.scala 51:27]
  reg [31:0] _RAND_320;
  reg  _T_996_1; // @[pearray.scala 51:27]
  reg [31:0] _RAND_321;
  reg  _T_996_2; // @[pearray.scala 51:27]
  reg [31:0] _RAND_322;
  reg  _T_996_3; // @[pearray.scala 51:27]
  reg [31:0] _RAND_323;
  reg  _T_1008_0; // @[pearray.scala 51:27]
  reg [31:0] _RAND_324;
  reg  _T_1008_1; // @[pearray.scala 51:27]
  reg [31:0] _RAND_325;
  reg  _T_1008_2; // @[pearray.scala 51:27]
  reg [31:0] _RAND_326;
  reg  _T_1008_3; // @[pearray.scala 51:27]
  reg [31:0] _RAND_327;
  reg  _T_1020_0; // @[pearray.scala 51:27]
  reg [31:0] _RAND_328;
  reg  _T_1020_1; // @[pearray.scala 51:27]
  reg [31:0] _RAND_329;
  reg  _T_1020_2; // @[pearray.scala 51:27]
  reg [31:0] _RAND_330;
  reg  _T_1020_3; // @[pearray.scala 51:27]
  reg [31:0] _RAND_331;
  reg  _T_1032_0; // @[pearray.scala 51:27]
  reg [31:0] _RAND_332;
  reg  _T_1032_1; // @[pearray.scala 51:27]
  reg [31:0] _RAND_333;
  reg  _T_1032_2; // @[pearray.scala 51:27]
  reg [31:0] _RAND_334;
  reg  _T_1032_3; // @[pearray.scala 51:27]
  reg [31:0] _RAND_335;
  reg  _T_1044_0; // @[pearray.scala 51:27]
  reg [31:0] _RAND_336;
  reg  _T_1044_1; // @[pearray.scala 51:27]
  reg [31:0] _RAND_337;
  reg  _T_1044_2; // @[pearray.scala 51:27]
  reg [31:0] _RAND_338;
  reg  _T_1044_3; // @[pearray.scala 51:27]
  reg [31:0] _RAND_339;
  reg  _T_1056_0; // @[pearray.scala 51:27]
  reg [31:0] _RAND_340;
  reg  _T_1056_1; // @[pearray.scala 51:27]
  reg [31:0] _RAND_341;
  reg  _T_1056_2; // @[pearray.scala 51:27]
  reg [31:0] _RAND_342;
  reg  _T_1056_3; // @[pearray.scala 51:27]
  reg [31:0] _RAND_343;
  reg  _T_1068_0; // @[pearray.scala 51:27]
  reg [31:0] _RAND_344;
  reg  _T_1068_1; // @[pearray.scala 51:27]
  reg [31:0] _RAND_345;
  reg  _T_1068_2; // @[pearray.scala 51:27]
  reg [31:0] _RAND_346;
  reg  _T_1068_3; // @[pearray.scala 51:27]
  reg [31:0] _RAND_347;
  wire  _T_1071 = MultiDimTime_io_index_1 == 18'h11; // @[pearray.scala 180:73]
  wire  _T_1073 = _T_1071 & _T_8; // @[pearray.scala 180:99]
  reg  _T_1080_0; // @[pearray.scala 51:27]
  reg [31:0] _RAND_348;
  reg  _T_1080_1; // @[pearray.scala 51:27]
  reg [31:0] _RAND_349;
  reg  _T_1080_2; // @[pearray.scala 51:27]
  reg [31:0] _RAND_350;
  reg  _T_1080_3; // @[pearray.scala 51:27]
  reg [31:0] _RAND_351;
  reg  _T_1094_0; // @[pearray.scala 51:27]
  reg [31:0] _RAND_352;
  reg  _T_1094_1; // @[pearray.scala 51:27]
  reg [31:0] _RAND_353;
  reg  _T_1094_2; // @[pearray.scala 51:27]
  reg [31:0] _RAND_354;
  reg  _T_1094_3; // @[pearray.scala 51:27]
  reg [31:0] _RAND_355;
  reg  _T_1106_0; // @[pearray.scala 51:27]
  reg [31:0] _RAND_356;
  reg  _T_1106_1; // @[pearray.scala 51:27]
  reg [31:0] _RAND_357;
  reg  _T_1106_2; // @[pearray.scala 51:27]
  reg [31:0] _RAND_358;
  reg  _T_1106_3; // @[pearray.scala 51:27]
  reg [31:0] _RAND_359;
  reg  _T_1118_0; // @[pearray.scala 51:27]
  reg [31:0] _RAND_360;
  reg  _T_1118_1; // @[pearray.scala 51:27]
  reg [31:0] _RAND_361;
  reg  _T_1118_2; // @[pearray.scala 51:27]
  reg [31:0] _RAND_362;
  reg  _T_1118_3; // @[pearray.scala 51:27]
  reg [31:0] _RAND_363;
  reg  _T_1130_0; // @[pearray.scala 51:27]
  reg [31:0] _RAND_364;
  reg  _T_1130_1; // @[pearray.scala 51:27]
  reg [31:0] _RAND_365;
  reg  _T_1130_2; // @[pearray.scala 51:27]
  reg [31:0] _RAND_366;
  reg  _T_1130_3; // @[pearray.scala 51:27]
  reg [31:0] _RAND_367;
  reg  _T_1142_0; // @[pearray.scala 51:27]
  reg [31:0] _RAND_368;
  reg  _T_1142_1; // @[pearray.scala 51:27]
  reg [31:0] _RAND_369;
  reg  _T_1142_2; // @[pearray.scala 51:27]
  reg [31:0] _RAND_370;
  reg  _T_1142_3; // @[pearray.scala 51:27]
  reg [31:0] _RAND_371;
  reg  _T_1154_0; // @[pearray.scala 51:27]
  reg [31:0] _RAND_372;
  reg  _T_1154_1; // @[pearray.scala 51:27]
  reg [31:0] _RAND_373;
  reg  _T_1154_2; // @[pearray.scala 51:27]
  reg [31:0] _RAND_374;
  reg  _T_1154_3; // @[pearray.scala 51:27]
  reg [31:0] _RAND_375;
  reg  _T_1166_0; // @[pearray.scala 51:27]
  reg [31:0] _RAND_376;
  reg  _T_1166_1; // @[pearray.scala 51:27]
  reg [31:0] _RAND_377;
  reg  _T_1166_2; // @[pearray.scala 51:27]
  reg [31:0] _RAND_378;
  reg  _T_1166_3; // @[pearray.scala 51:27]
  reg [31:0] _RAND_379;
  wire  _T_1169 = MultiDimTime_io_index_1 == 18'h12; // @[pearray.scala 180:73]
  wire  _T_1171 = _T_1169 & _T_8; // @[pearray.scala 180:99]
  reg  _T_1178_0; // @[pearray.scala 51:27]
  reg [31:0] _RAND_380;
  reg  _T_1178_1; // @[pearray.scala 51:27]
  reg [31:0] _RAND_381;
  reg  _T_1178_2; // @[pearray.scala 51:27]
  reg [31:0] _RAND_382;
  reg  _T_1178_3; // @[pearray.scala 51:27]
  reg [31:0] _RAND_383;
  reg  _T_1192_0; // @[pearray.scala 51:27]
  reg [31:0] _RAND_384;
  reg  _T_1192_1; // @[pearray.scala 51:27]
  reg [31:0] _RAND_385;
  reg  _T_1192_2; // @[pearray.scala 51:27]
  reg [31:0] _RAND_386;
  reg  _T_1192_3; // @[pearray.scala 51:27]
  reg [31:0] _RAND_387;
  reg  _T_1204_0; // @[pearray.scala 51:27]
  reg [31:0] _RAND_388;
  reg  _T_1204_1; // @[pearray.scala 51:27]
  reg [31:0] _RAND_389;
  reg  _T_1204_2; // @[pearray.scala 51:27]
  reg [31:0] _RAND_390;
  reg  _T_1204_3; // @[pearray.scala 51:27]
  reg [31:0] _RAND_391;
  reg  _T_1216_0; // @[pearray.scala 51:27]
  reg [31:0] _RAND_392;
  reg  _T_1216_1; // @[pearray.scala 51:27]
  reg [31:0] _RAND_393;
  reg  _T_1216_2; // @[pearray.scala 51:27]
  reg [31:0] _RAND_394;
  reg  _T_1216_3; // @[pearray.scala 51:27]
  reg [31:0] _RAND_395;
  reg  _T_1228_0; // @[pearray.scala 51:27]
  reg [31:0] _RAND_396;
  reg  _T_1228_1; // @[pearray.scala 51:27]
  reg [31:0] _RAND_397;
  reg  _T_1228_2; // @[pearray.scala 51:27]
  reg [31:0] _RAND_398;
  reg  _T_1228_3; // @[pearray.scala 51:27]
  reg [31:0] _RAND_399;
  reg  _T_1240_0; // @[pearray.scala 51:27]
  reg [31:0] _RAND_400;
  reg  _T_1240_1; // @[pearray.scala 51:27]
  reg [31:0] _RAND_401;
  reg  _T_1240_2; // @[pearray.scala 51:27]
  reg [31:0] _RAND_402;
  reg  _T_1240_3; // @[pearray.scala 51:27]
  reg [31:0] _RAND_403;
  reg  _T_1252_0; // @[pearray.scala 51:27]
  reg [31:0] _RAND_404;
  reg  _T_1252_1; // @[pearray.scala 51:27]
  reg [31:0] _RAND_405;
  reg  _T_1252_2; // @[pearray.scala 51:27]
  reg [31:0] _RAND_406;
  reg  _T_1252_3; // @[pearray.scala 51:27]
  reg [31:0] _RAND_407;
  reg  _T_1264_0; // @[pearray.scala 51:27]
  reg [31:0] _RAND_408;
  reg  _T_1264_1; // @[pearray.scala 51:27]
  reg [31:0] _RAND_409;
  reg  _T_1264_2; // @[pearray.scala 51:27]
  reg [31:0] _RAND_410;
  reg  _T_1264_3; // @[pearray.scala 51:27]
  reg [31:0] _RAND_411;
  wire  _T_1267 = MultiDimTime_io_index_1 == 18'h13; // @[pearray.scala 180:73]
  wire  _T_1269 = _T_1267 & _T_8; // @[pearray.scala 180:99]
  reg  _T_1276_0; // @[pearray.scala 51:27]
  reg [31:0] _RAND_412;
  reg  _T_1276_1; // @[pearray.scala 51:27]
  reg [31:0] _RAND_413;
  reg  _T_1276_2; // @[pearray.scala 51:27]
  reg [31:0] _RAND_414;
  reg  _T_1276_3; // @[pearray.scala 51:27]
  reg [31:0] _RAND_415;
  reg  _T_1290_0; // @[pearray.scala 51:27]
  reg [31:0] _RAND_416;
  reg  _T_1290_1; // @[pearray.scala 51:27]
  reg [31:0] _RAND_417;
  reg  _T_1290_2; // @[pearray.scala 51:27]
  reg [31:0] _RAND_418;
  reg  _T_1290_3; // @[pearray.scala 51:27]
  reg [31:0] _RAND_419;
  reg  _T_1302_0; // @[pearray.scala 51:27]
  reg [31:0] _RAND_420;
  reg  _T_1302_1; // @[pearray.scala 51:27]
  reg [31:0] _RAND_421;
  reg  _T_1302_2; // @[pearray.scala 51:27]
  reg [31:0] _RAND_422;
  reg  _T_1302_3; // @[pearray.scala 51:27]
  reg [31:0] _RAND_423;
  reg  _T_1314_0; // @[pearray.scala 51:27]
  reg [31:0] _RAND_424;
  reg  _T_1314_1; // @[pearray.scala 51:27]
  reg [31:0] _RAND_425;
  reg  _T_1314_2; // @[pearray.scala 51:27]
  reg [31:0] _RAND_426;
  reg  _T_1314_3; // @[pearray.scala 51:27]
  reg [31:0] _RAND_427;
  reg  _T_1326_0; // @[pearray.scala 51:27]
  reg [31:0] _RAND_428;
  reg  _T_1326_1; // @[pearray.scala 51:27]
  reg [31:0] _RAND_429;
  reg  _T_1326_2; // @[pearray.scala 51:27]
  reg [31:0] _RAND_430;
  reg  _T_1326_3; // @[pearray.scala 51:27]
  reg [31:0] _RAND_431;
  reg  _T_1338_0; // @[pearray.scala 51:27]
  reg [31:0] _RAND_432;
  reg  _T_1338_1; // @[pearray.scala 51:27]
  reg [31:0] _RAND_433;
  reg  _T_1338_2; // @[pearray.scala 51:27]
  reg [31:0] _RAND_434;
  reg  _T_1338_3; // @[pearray.scala 51:27]
  reg [31:0] _RAND_435;
  reg  _T_1350_0; // @[pearray.scala 51:27]
  reg [31:0] _RAND_436;
  reg  _T_1350_1; // @[pearray.scala 51:27]
  reg [31:0] _RAND_437;
  reg  _T_1350_2; // @[pearray.scala 51:27]
  reg [31:0] _RAND_438;
  reg  _T_1350_3; // @[pearray.scala 51:27]
  reg [31:0] _RAND_439;
  reg  _T_1362_0; // @[pearray.scala 51:27]
  reg [31:0] _RAND_440;
  reg  _T_1362_1; // @[pearray.scala 51:27]
  reg [31:0] _RAND_441;
  reg  _T_1362_2; // @[pearray.scala 51:27]
  reg [31:0] _RAND_442;
  reg  _T_1362_3; // @[pearray.scala 51:27]
  reg [31:0] _RAND_443;
  wire  _T_1365 = MultiDimTime_io_index_1 == 18'h14; // @[pearray.scala 180:73]
  wire  _T_1367 = _T_1365 & _T_8; // @[pearray.scala 180:99]
  reg  _T_1374_0; // @[pearray.scala 51:27]
  reg [31:0] _RAND_444;
  reg  _T_1374_1; // @[pearray.scala 51:27]
  reg [31:0] _RAND_445;
  reg  _T_1374_2; // @[pearray.scala 51:27]
  reg [31:0] _RAND_446;
  reg  _T_1374_3; // @[pearray.scala 51:27]
  reg [31:0] _RAND_447;
  reg  _T_1388_0; // @[pearray.scala 51:27]
  reg [31:0] _RAND_448;
  reg  _T_1388_1; // @[pearray.scala 51:27]
  reg [31:0] _RAND_449;
  reg  _T_1388_2; // @[pearray.scala 51:27]
  reg [31:0] _RAND_450;
  reg  _T_1388_3; // @[pearray.scala 51:27]
  reg [31:0] _RAND_451;
  reg  _T_1400_0; // @[pearray.scala 51:27]
  reg [31:0] _RAND_452;
  reg  _T_1400_1; // @[pearray.scala 51:27]
  reg [31:0] _RAND_453;
  reg  _T_1400_2; // @[pearray.scala 51:27]
  reg [31:0] _RAND_454;
  reg  _T_1400_3; // @[pearray.scala 51:27]
  reg [31:0] _RAND_455;
  reg  _T_1412_0; // @[pearray.scala 51:27]
  reg [31:0] _RAND_456;
  reg  _T_1412_1; // @[pearray.scala 51:27]
  reg [31:0] _RAND_457;
  reg  _T_1412_2; // @[pearray.scala 51:27]
  reg [31:0] _RAND_458;
  reg  _T_1412_3; // @[pearray.scala 51:27]
  reg [31:0] _RAND_459;
  reg  _T_1424_0; // @[pearray.scala 51:27]
  reg [31:0] _RAND_460;
  reg  _T_1424_1; // @[pearray.scala 51:27]
  reg [31:0] _RAND_461;
  reg  _T_1424_2; // @[pearray.scala 51:27]
  reg [31:0] _RAND_462;
  reg  _T_1424_3; // @[pearray.scala 51:27]
  reg [31:0] _RAND_463;
  reg  _T_1436_0; // @[pearray.scala 51:27]
  reg [31:0] _RAND_464;
  reg  _T_1436_1; // @[pearray.scala 51:27]
  reg [31:0] _RAND_465;
  reg  _T_1436_2; // @[pearray.scala 51:27]
  reg [31:0] _RAND_466;
  reg  _T_1436_3; // @[pearray.scala 51:27]
  reg [31:0] _RAND_467;
  reg  _T_1448_0; // @[pearray.scala 51:27]
  reg [31:0] _RAND_468;
  reg  _T_1448_1; // @[pearray.scala 51:27]
  reg [31:0] _RAND_469;
  reg  _T_1448_2; // @[pearray.scala 51:27]
  reg [31:0] _RAND_470;
  reg  _T_1448_3; // @[pearray.scala 51:27]
  reg [31:0] _RAND_471;
  reg  _T_1460_0; // @[pearray.scala 51:27]
  reg [31:0] _RAND_472;
  reg  _T_1460_1; // @[pearray.scala 51:27]
  reg [31:0] _RAND_473;
  reg  _T_1460_2; // @[pearray.scala 51:27]
  reg [31:0] _RAND_474;
  reg  _T_1460_3; // @[pearray.scala 51:27]
  reg [31:0] _RAND_475;
  wire  _T_1463 = MultiDimTime_io_index_1 == 18'h15; // @[pearray.scala 180:73]
  wire  _T_1465 = _T_1463 & _T_8; // @[pearray.scala 180:99]
  reg  _T_1472_0; // @[pearray.scala 51:27]
  reg [31:0] _RAND_476;
  reg  _T_1472_1; // @[pearray.scala 51:27]
  reg [31:0] _RAND_477;
  reg  _T_1472_2; // @[pearray.scala 51:27]
  reg [31:0] _RAND_478;
  reg  _T_1472_3; // @[pearray.scala 51:27]
  reg [31:0] _RAND_479;
  reg  _T_1486_0; // @[pearray.scala 51:27]
  reg [31:0] _RAND_480;
  reg  _T_1486_1; // @[pearray.scala 51:27]
  reg [31:0] _RAND_481;
  reg  _T_1486_2; // @[pearray.scala 51:27]
  reg [31:0] _RAND_482;
  reg  _T_1486_3; // @[pearray.scala 51:27]
  reg [31:0] _RAND_483;
  reg  _T_1498_0; // @[pearray.scala 51:27]
  reg [31:0] _RAND_484;
  reg  _T_1498_1; // @[pearray.scala 51:27]
  reg [31:0] _RAND_485;
  reg  _T_1498_2; // @[pearray.scala 51:27]
  reg [31:0] _RAND_486;
  reg  _T_1498_3; // @[pearray.scala 51:27]
  reg [31:0] _RAND_487;
  reg  _T_1510_0; // @[pearray.scala 51:27]
  reg [31:0] _RAND_488;
  reg  _T_1510_1; // @[pearray.scala 51:27]
  reg [31:0] _RAND_489;
  reg  _T_1510_2; // @[pearray.scala 51:27]
  reg [31:0] _RAND_490;
  reg  _T_1510_3; // @[pearray.scala 51:27]
  reg [31:0] _RAND_491;
  reg  _T_1522_0; // @[pearray.scala 51:27]
  reg [31:0] _RAND_492;
  reg  _T_1522_1; // @[pearray.scala 51:27]
  reg [31:0] _RAND_493;
  reg  _T_1522_2; // @[pearray.scala 51:27]
  reg [31:0] _RAND_494;
  reg  _T_1522_3; // @[pearray.scala 51:27]
  reg [31:0] _RAND_495;
  reg  _T_1534_0; // @[pearray.scala 51:27]
  reg [31:0] _RAND_496;
  reg  _T_1534_1; // @[pearray.scala 51:27]
  reg [31:0] _RAND_497;
  reg  _T_1534_2; // @[pearray.scala 51:27]
  reg [31:0] _RAND_498;
  reg  _T_1534_3; // @[pearray.scala 51:27]
  reg [31:0] _RAND_499;
  reg  _T_1546_0; // @[pearray.scala 51:27]
  reg [31:0] _RAND_500;
  reg  _T_1546_1; // @[pearray.scala 51:27]
  reg [31:0] _RAND_501;
  reg  _T_1546_2; // @[pearray.scala 51:27]
  reg [31:0] _RAND_502;
  reg  _T_1546_3; // @[pearray.scala 51:27]
  reg [31:0] _RAND_503;
  reg  _T_1558_0; // @[pearray.scala 51:27]
  reg [31:0] _RAND_504;
  reg  _T_1558_1; // @[pearray.scala 51:27]
  reg [31:0] _RAND_505;
  reg  _T_1558_2; // @[pearray.scala 51:27]
  reg [31:0] _RAND_506;
  reg  _T_1558_3; // @[pearray.scala 51:27]
  reg [31:0] _RAND_507;
  wire  _T_1561 = MultiDimTime_io_index_1 == 18'h16; // @[pearray.scala 180:73]
  wire  _T_1563 = _T_1561 & _T_8; // @[pearray.scala 180:99]
  reg  _T_1570_0; // @[pearray.scala 51:27]
  reg [31:0] _RAND_508;
  reg  _T_1570_1; // @[pearray.scala 51:27]
  reg [31:0] _RAND_509;
  reg  _T_1570_2; // @[pearray.scala 51:27]
  reg [31:0] _RAND_510;
  reg  _T_1570_3; // @[pearray.scala 51:27]
  reg [31:0] _RAND_511;
  wire  _T_1579 = MultiDimTime_io_index_1 < 18'h8; // @[pearray.scala 236:134]
  wire  _T_1580 = io_exec_valid & _T_1579; // @[pearray.scala 236:112]
  reg  _T_1585_0; // @[pearray.scala 51:27]
  reg [31:0] _RAND_512;
  reg  _T_1585_1; // @[pearray.scala 51:27]
  reg [31:0] _RAND_513;
  reg  _T_1585_2; // @[pearray.scala 51:27]
  reg [31:0] _RAND_514;
  wire  _T_1586 = MultiDimTime_io_index_1 >= 18'h1; // @[pearray.scala 236:82]
  wire  _T_1587 = io_exec_valid & _T_1586; // @[pearray.scala 236:60]
  wire  _T_1588 = MultiDimTime_io_index_1 < 18'h9; // @[pearray.scala 236:134]
  wire  _T_1589 = _T_1587 & _T_1588; // @[pearray.scala 236:112]
  reg  _T_1594_0; // @[pearray.scala 51:27]
  reg [31:0] _RAND_515;
  reg  _T_1594_1; // @[pearray.scala 51:27]
  reg [31:0] _RAND_516;
  reg  _T_1594_2; // @[pearray.scala 51:27]
  reg [31:0] _RAND_517;
  wire  _T_1595 = MultiDimTime_io_index_1 >= 18'h2; // @[pearray.scala 236:82]
  wire  _T_1596 = io_exec_valid & _T_1595; // @[pearray.scala 236:60]
  wire  _T_1597 = MultiDimTime_io_index_1 < 18'ha; // @[pearray.scala 236:134]
  wire  _T_1598 = _T_1596 & _T_1597; // @[pearray.scala 236:112]
  reg  _T_1603_0; // @[pearray.scala 51:27]
  reg [31:0] _RAND_518;
  reg  _T_1603_1; // @[pearray.scala 51:27]
  reg [31:0] _RAND_519;
  reg  _T_1603_2; // @[pearray.scala 51:27]
  reg [31:0] _RAND_520;
  wire  _T_1604 = MultiDimTime_io_index_1 >= 18'h3; // @[pearray.scala 236:82]
  wire  _T_1605 = io_exec_valid & _T_1604; // @[pearray.scala 236:60]
  wire  _T_1606 = MultiDimTime_io_index_1 < 18'hb; // @[pearray.scala 236:134]
  wire  _T_1607 = _T_1605 & _T_1606; // @[pearray.scala 236:112]
  reg  _T_1612_0; // @[pearray.scala 51:27]
  reg [31:0] _RAND_521;
  reg  _T_1612_1; // @[pearray.scala 51:27]
  reg [31:0] _RAND_522;
  reg  _T_1612_2; // @[pearray.scala 51:27]
  reg [31:0] _RAND_523;
  wire  _T_1613 = MultiDimTime_io_index_1 >= 18'h4; // @[pearray.scala 236:82]
  wire  _T_1614 = io_exec_valid & _T_1613; // @[pearray.scala 236:60]
  wire  _T_1615 = MultiDimTime_io_index_1 < 18'hc; // @[pearray.scala 236:134]
  wire  _T_1616 = _T_1614 & _T_1615; // @[pearray.scala 236:112]
  reg  _T_1621_0; // @[pearray.scala 51:27]
  reg [31:0] _RAND_524;
  reg  _T_1621_1; // @[pearray.scala 51:27]
  reg [31:0] _RAND_525;
  reg  _T_1621_2; // @[pearray.scala 51:27]
  reg [31:0] _RAND_526;
  wire  _T_1622 = MultiDimTime_io_index_1 >= 18'h5; // @[pearray.scala 236:82]
  wire  _T_1623 = io_exec_valid & _T_1622; // @[pearray.scala 236:60]
  wire  _T_1624 = MultiDimTime_io_index_1 < 18'hd; // @[pearray.scala 236:134]
  wire  _T_1625 = _T_1623 & _T_1624; // @[pearray.scala 236:112]
  reg  _T_1630_0; // @[pearray.scala 51:27]
  reg [31:0] _RAND_527;
  reg  _T_1630_1; // @[pearray.scala 51:27]
  reg [31:0] _RAND_528;
  reg  _T_1630_2; // @[pearray.scala 51:27]
  reg [31:0] _RAND_529;
  wire  _T_1631 = MultiDimTime_io_index_1 >= 18'h6; // @[pearray.scala 236:82]
  wire  _T_1632 = io_exec_valid & _T_1631; // @[pearray.scala 236:60]
  wire  _T_1633 = MultiDimTime_io_index_1 < 18'he; // @[pearray.scala 236:134]
  wire  _T_1634 = _T_1632 & _T_1633; // @[pearray.scala 236:112]
  reg  _T_1639_0; // @[pearray.scala 51:27]
  reg [31:0] _RAND_530;
  reg  _T_1639_1; // @[pearray.scala 51:27]
  reg [31:0] _RAND_531;
  reg  _T_1639_2; // @[pearray.scala 51:27]
  reg [31:0] _RAND_532;
  wire  _T_1640 = MultiDimTime_io_index_1 >= 18'h7; // @[pearray.scala 236:82]
  wire  _T_1641 = io_exec_valid & _T_1640; // @[pearray.scala 236:60]
  wire  _T_1642 = MultiDimTime_io_index_1 < 18'hf; // @[pearray.scala 236:134]
  wire  _T_1643 = _T_1641 & _T_1642; // @[pearray.scala 236:112]
  reg  _T_1648_0; // @[pearray.scala 51:27]
  reg [31:0] _RAND_533;
  reg  _T_1648_1; // @[pearray.scala 51:27]
  reg [31:0] _RAND_534;
  reg  _T_1648_2; // @[pearray.scala 51:27]
  reg [31:0] _RAND_535;
  wire  _T_1649 = MultiDimTime_io_index_1 >= 18'h8; // @[pearray.scala 236:82]
  wire  _T_1650 = io_exec_valid & _T_1649; // @[pearray.scala 236:60]
  wire  _T_1651 = MultiDimTime_io_index_1 < 18'h10; // @[pearray.scala 236:134]
  wire  _T_1652 = _T_1650 & _T_1651; // @[pearray.scala 236:112]
  reg  _T_1657_0; // @[pearray.scala 51:27]
  reg [31:0] _RAND_536;
  reg  _T_1657_1; // @[pearray.scala 51:27]
  reg [31:0] _RAND_537;
  reg  _T_1657_2; // @[pearray.scala 51:27]
  reg [31:0] _RAND_538;
  wire  _T_1658 = MultiDimTime_io_index_1 >= 18'h9; // @[pearray.scala 236:82]
  wire  _T_1659 = io_exec_valid & _T_1658; // @[pearray.scala 236:60]
  wire  _T_1660 = MultiDimTime_io_index_1 < 18'h11; // @[pearray.scala 236:134]
  wire  _T_1661 = _T_1659 & _T_1660; // @[pearray.scala 236:112]
  reg  _T_1666_0; // @[pearray.scala 51:27]
  reg [31:0] _RAND_539;
  reg  _T_1666_1; // @[pearray.scala 51:27]
  reg [31:0] _RAND_540;
  reg  _T_1666_2; // @[pearray.scala 51:27]
  reg [31:0] _RAND_541;
  wire  _T_1667 = MultiDimTime_io_index_1 >= 18'ha; // @[pearray.scala 236:82]
  wire  _T_1668 = io_exec_valid & _T_1667; // @[pearray.scala 236:60]
  wire  _T_1669 = MultiDimTime_io_index_1 < 18'h12; // @[pearray.scala 236:134]
  wire  _T_1670 = _T_1668 & _T_1669; // @[pearray.scala 236:112]
  reg  _T_1675_0; // @[pearray.scala 51:27]
  reg [31:0] _RAND_542;
  reg  _T_1675_1; // @[pearray.scala 51:27]
  reg [31:0] _RAND_543;
  reg  _T_1675_2; // @[pearray.scala 51:27]
  reg [31:0] _RAND_544;
  wire  _T_1676 = MultiDimTime_io_index_1 >= 18'hb; // @[pearray.scala 236:82]
  wire  _T_1677 = io_exec_valid & _T_1676; // @[pearray.scala 236:60]
  wire  _T_1678 = MultiDimTime_io_index_1 < 18'h13; // @[pearray.scala 236:134]
  wire  _T_1679 = _T_1677 & _T_1678; // @[pearray.scala 236:112]
  reg  _T_1684_0; // @[pearray.scala 51:27]
  reg [31:0] _RAND_545;
  reg  _T_1684_1; // @[pearray.scala 51:27]
  reg [31:0] _RAND_546;
  reg  _T_1684_2; // @[pearray.scala 51:27]
  reg [31:0] _RAND_547;
  wire  _T_1685 = MultiDimTime_io_index_1 >= 18'hc; // @[pearray.scala 236:82]
  wire  _T_1686 = io_exec_valid & _T_1685; // @[pearray.scala 236:60]
  wire  _T_1687 = MultiDimTime_io_index_1 < 18'h14; // @[pearray.scala 236:134]
  wire  _T_1688 = _T_1686 & _T_1687; // @[pearray.scala 236:112]
  reg  _T_1693_0; // @[pearray.scala 51:27]
  reg [31:0] _RAND_548;
  reg  _T_1693_1; // @[pearray.scala 51:27]
  reg [31:0] _RAND_549;
  reg  _T_1693_2; // @[pearray.scala 51:27]
  reg [31:0] _RAND_550;
  wire  _T_1694 = MultiDimTime_io_index_1 >= 18'hd; // @[pearray.scala 236:82]
  wire  _T_1695 = io_exec_valid & _T_1694; // @[pearray.scala 236:60]
  wire  _T_1696 = MultiDimTime_io_index_1 < 18'h15; // @[pearray.scala 236:134]
  wire  _T_1697 = _T_1695 & _T_1696; // @[pearray.scala 236:112]
  reg  _T_1702_0; // @[pearray.scala 51:27]
  reg [31:0] _RAND_551;
  reg  _T_1702_1; // @[pearray.scala 51:27]
  reg [31:0] _RAND_552;
  reg  _T_1702_2; // @[pearray.scala 51:27]
  reg [31:0] _RAND_553;
  wire  _T_1703 = MultiDimTime_io_index_1 >= 18'he; // @[pearray.scala 236:82]
  wire  _T_1704 = io_exec_valid & _T_1703; // @[pearray.scala 236:60]
  wire  _T_1705 = MultiDimTime_io_index_1 < 18'h16; // @[pearray.scala 236:134]
  wire  _T_1706 = _T_1704 & _T_1705; // @[pearray.scala 236:112]
  reg  _T_1711_0; // @[pearray.scala 51:27]
  reg [31:0] _RAND_554;
  reg  _T_1711_1; // @[pearray.scala 51:27]
  reg [31:0] _RAND_555;
  reg  _T_1711_2; // @[pearray.scala 51:27]
  reg [31:0] _RAND_556;
  wire  _T_1712 = MultiDimTime_io_index_1 >= 18'hf; // @[pearray.scala 236:82]
  wire  _T_1713 = io_exec_valid & _T_1712; // @[pearray.scala 236:60]
  wire  _T_1714 = MultiDimTime_io_index_1 < 18'h17; // @[pearray.scala 236:134]
  wire  _T_1715 = _T_1713 & _T_1714; // @[pearray.scala 236:112]
  reg  _T_1720_0; // @[pearray.scala 51:27]
  reg [31:0] _RAND_557;
  reg  _T_1720_1; // @[pearray.scala 51:27]
  reg [31:0] _RAND_558;
  reg  _T_1720_2; // @[pearray.scala 51:27]
  reg [31:0] _RAND_559;
  reg  _T_1722_0; // @[pearray.scala 213:27]
  reg [31:0] _RAND_560;
  reg  _T_1722_1; // @[pearray.scala 213:27]
  reg [31:0] _RAND_561;
  reg  _T_1722_2; // @[pearray.scala 213:27]
  reg [31:0] _RAND_562;
  reg  _T_1722_3; // @[pearray.scala 213:27]
  reg [31:0] _RAND_563;
  reg  _T_1722_4; // @[pearray.scala 213:27]
  reg [31:0] _RAND_564;
  reg  _T_1722_5; // @[pearray.scala 213:27]
  reg [31:0] _RAND_565;
  reg  _T_1722_6; // @[pearray.scala 213:27]
  reg [31:0] _RAND_566;
  MultiDimTime MultiDimTime ( // @[pearray.scala 63:25]
    .clock(MultiDimTime_clock),
    .reset(MultiDimTime_reset),
    .io_in(MultiDimTime_io_in),
    .io_out_0(MultiDimTime_io_out_0),
    .io_out_1(MultiDimTime_io_out_1),
    .io_index_0(MultiDimTime_io_index_0),
    .io_index_1(MultiDimTime_io_index_1)
  );
  PE PE ( // @[pearray.scala 101:13]
    .clock(PE_clock),
    .reset(PE_reset),
    .io_data_2_in_bits(PE_io_data_2_in_bits),
    .io_data_2_out_bits(PE_io_data_2_out_bits),
    .io_data_1_in_valid(PE_io_data_1_in_valid),
    .io_data_1_in_bits(PE_io_data_1_in_bits),
    .io_data_1_out_valid(PE_io_data_1_out_valid),
    .io_data_1_out_bits(PE_io_data_1_out_bits),
    .io_data_0_in_valid(PE_io_data_0_in_valid),
    .io_data_0_in_bits(PE_io_data_0_in_bits),
    .io_data_0_out_valid(PE_io_data_0_out_valid),
    .io_data_0_out_bits(PE_io_data_0_out_bits),
    .io_sig_stat2trans(PE_io_sig_stat2trans)
  );
  PE PE_1 ( // @[pearray.scala 101:13]
    .clock(PE_1_clock),
    .reset(PE_1_reset),
    .io_data_2_in_bits(PE_1_io_data_2_in_bits),
    .io_data_2_out_bits(PE_1_io_data_2_out_bits),
    .io_data_1_in_valid(PE_1_io_data_1_in_valid),
    .io_data_1_in_bits(PE_1_io_data_1_in_bits),
    .io_data_1_out_valid(PE_1_io_data_1_out_valid),
    .io_data_1_out_bits(PE_1_io_data_1_out_bits),
    .io_data_0_in_valid(PE_1_io_data_0_in_valid),
    .io_data_0_in_bits(PE_1_io_data_0_in_bits),
    .io_data_0_out_valid(PE_1_io_data_0_out_valid),
    .io_data_0_out_bits(PE_1_io_data_0_out_bits),
    .io_sig_stat2trans(PE_1_io_sig_stat2trans)
  );
  PE PE_2 ( // @[pearray.scala 101:13]
    .clock(PE_2_clock),
    .reset(PE_2_reset),
    .io_data_2_in_bits(PE_2_io_data_2_in_bits),
    .io_data_2_out_bits(PE_2_io_data_2_out_bits),
    .io_data_1_in_valid(PE_2_io_data_1_in_valid),
    .io_data_1_in_bits(PE_2_io_data_1_in_bits),
    .io_data_1_out_valid(PE_2_io_data_1_out_valid),
    .io_data_1_out_bits(PE_2_io_data_1_out_bits),
    .io_data_0_in_valid(PE_2_io_data_0_in_valid),
    .io_data_0_in_bits(PE_2_io_data_0_in_bits),
    .io_data_0_out_valid(PE_2_io_data_0_out_valid),
    .io_data_0_out_bits(PE_2_io_data_0_out_bits),
    .io_sig_stat2trans(PE_2_io_sig_stat2trans)
  );
  PE PE_3 ( // @[pearray.scala 101:13]
    .clock(PE_3_clock),
    .reset(PE_3_reset),
    .io_data_2_in_bits(PE_3_io_data_2_in_bits),
    .io_data_2_out_bits(PE_3_io_data_2_out_bits),
    .io_data_1_in_valid(PE_3_io_data_1_in_valid),
    .io_data_1_in_bits(PE_3_io_data_1_in_bits),
    .io_data_1_out_valid(PE_3_io_data_1_out_valid),
    .io_data_1_out_bits(PE_3_io_data_1_out_bits),
    .io_data_0_in_valid(PE_3_io_data_0_in_valid),
    .io_data_0_in_bits(PE_3_io_data_0_in_bits),
    .io_data_0_out_valid(PE_3_io_data_0_out_valid),
    .io_data_0_out_bits(PE_3_io_data_0_out_bits),
    .io_sig_stat2trans(PE_3_io_sig_stat2trans)
  );
  PE PE_4 ( // @[pearray.scala 101:13]
    .clock(PE_4_clock),
    .reset(PE_4_reset),
    .io_data_2_in_bits(PE_4_io_data_2_in_bits),
    .io_data_2_out_bits(PE_4_io_data_2_out_bits),
    .io_data_1_in_valid(PE_4_io_data_1_in_valid),
    .io_data_1_in_bits(PE_4_io_data_1_in_bits),
    .io_data_1_out_valid(PE_4_io_data_1_out_valid),
    .io_data_1_out_bits(PE_4_io_data_1_out_bits),
    .io_data_0_in_valid(PE_4_io_data_0_in_valid),
    .io_data_0_in_bits(PE_4_io_data_0_in_bits),
    .io_data_0_out_valid(PE_4_io_data_0_out_valid),
    .io_data_0_out_bits(PE_4_io_data_0_out_bits),
    .io_sig_stat2trans(PE_4_io_sig_stat2trans)
  );
  PE PE_5 ( // @[pearray.scala 101:13]
    .clock(PE_5_clock),
    .reset(PE_5_reset),
    .io_data_2_in_bits(PE_5_io_data_2_in_bits),
    .io_data_2_out_bits(PE_5_io_data_2_out_bits),
    .io_data_1_in_valid(PE_5_io_data_1_in_valid),
    .io_data_1_in_bits(PE_5_io_data_1_in_bits),
    .io_data_1_out_valid(PE_5_io_data_1_out_valid),
    .io_data_1_out_bits(PE_5_io_data_1_out_bits),
    .io_data_0_in_valid(PE_5_io_data_0_in_valid),
    .io_data_0_in_bits(PE_5_io_data_0_in_bits),
    .io_data_0_out_valid(PE_5_io_data_0_out_valid),
    .io_data_0_out_bits(PE_5_io_data_0_out_bits),
    .io_sig_stat2trans(PE_5_io_sig_stat2trans)
  );
  PE PE_6 ( // @[pearray.scala 101:13]
    .clock(PE_6_clock),
    .reset(PE_6_reset),
    .io_data_2_in_bits(PE_6_io_data_2_in_bits),
    .io_data_2_out_bits(PE_6_io_data_2_out_bits),
    .io_data_1_in_valid(PE_6_io_data_1_in_valid),
    .io_data_1_in_bits(PE_6_io_data_1_in_bits),
    .io_data_1_out_valid(PE_6_io_data_1_out_valid),
    .io_data_1_out_bits(PE_6_io_data_1_out_bits),
    .io_data_0_in_valid(PE_6_io_data_0_in_valid),
    .io_data_0_in_bits(PE_6_io_data_0_in_bits),
    .io_data_0_out_valid(PE_6_io_data_0_out_valid),
    .io_data_0_out_bits(PE_6_io_data_0_out_bits),
    .io_sig_stat2trans(PE_6_io_sig_stat2trans)
  );
  PE PE_7 ( // @[pearray.scala 101:13]
    .clock(PE_7_clock),
    .reset(PE_7_reset),
    .io_data_2_in_bits(PE_7_io_data_2_in_bits),
    .io_data_2_out_bits(PE_7_io_data_2_out_bits),
    .io_data_1_in_valid(PE_7_io_data_1_in_valid),
    .io_data_1_in_bits(PE_7_io_data_1_in_bits),
    .io_data_1_out_valid(PE_7_io_data_1_out_valid),
    .io_data_1_out_bits(PE_7_io_data_1_out_bits),
    .io_data_0_in_valid(PE_7_io_data_0_in_valid),
    .io_data_0_in_bits(PE_7_io_data_0_in_bits),
    .io_data_0_out_valid(PE_7_io_data_0_out_valid),
    .io_data_0_out_bits(PE_7_io_data_0_out_bits),
    .io_sig_stat2trans(PE_7_io_sig_stat2trans)
  );
  PE PE_8 ( // @[pearray.scala 101:13]
    .clock(PE_8_clock),
    .reset(PE_8_reset),
    .io_data_2_in_bits(PE_8_io_data_2_in_bits),
    .io_data_2_out_bits(PE_8_io_data_2_out_bits),
    .io_data_1_in_valid(PE_8_io_data_1_in_valid),
    .io_data_1_in_bits(PE_8_io_data_1_in_bits),
    .io_data_1_out_valid(PE_8_io_data_1_out_valid),
    .io_data_1_out_bits(PE_8_io_data_1_out_bits),
    .io_data_0_in_valid(PE_8_io_data_0_in_valid),
    .io_data_0_in_bits(PE_8_io_data_0_in_bits),
    .io_data_0_out_valid(PE_8_io_data_0_out_valid),
    .io_data_0_out_bits(PE_8_io_data_0_out_bits),
    .io_sig_stat2trans(PE_8_io_sig_stat2trans)
  );
  PE PE_9 ( // @[pearray.scala 101:13]
    .clock(PE_9_clock),
    .reset(PE_9_reset),
    .io_data_2_in_bits(PE_9_io_data_2_in_bits),
    .io_data_2_out_bits(PE_9_io_data_2_out_bits),
    .io_data_1_in_valid(PE_9_io_data_1_in_valid),
    .io_data_1_in_bits(PE_9_io_data_1_in_bits),
    .io_data_1_out_valid(PE_9_io_data_1_out_valid),
    .io_data_1_out_bits(PE_9_io_data_1_out_bits),
    .io_data_0_in_valid(PE_9_io_data_0_in_valid),
    .io_data_0_in_bits(PE_9_io_data_0_in_bits),
    .io_data_0_out_valid(PE_9_io_data_0_out_valid),
    .io_data_0_out_bits(PE_9_io_data_0_out_bits),
    .io_sig_stat2trans(PE_9_io_sig_stat2trans)
  );
  PE PE_10 ( // @[pearray.scala 101:13]
    .clock(PE_10_clock),
    .reset(PE_10_reset),
    .io_data_2_in_bits(PE_10_io_data_2_in_bits),
    .io_data_2_out_bits(PE_10_io_data_2_out_bits),
    .io_data_1_in_valid(PE_10_io_data_1_in_valid),
    .io_data_1_in_bits(PE_10_io_data_1_in_bits),
    .io_data_1_out_valid(PE_10_io_data_1_out_valid),
    .io_data_1_out_bits(PE_10_io_data_1_out_bits),
    .io_data_0_in_valid(PE_10_io_data_0_in_valid),
    .io_data_0_in_bits(PE_10_io_data_0_in_bits),
    .io_data_0_out_valid(PE_10_io_data_0_out_valid),
    .io_data_0_out_bits(PE_10_io_data_0_out_bits),
    .io_sig_stat2trans(PE_10_io_sig_stat2trans)
  );
  PE PE_11 ( // @[pearray.scala 101:13]
    .clock(PE_11_clock),
    .reset(PE_11_reset),
    .io_data_2_in_bits(PE_11_io_data_2_in_bits),
    .io_data_2_out_bits(PE_11_io_data_2_out_bits),
    .io_data_1_in_valid(PE_11_io_data_1_in_valid),
    .io_data_1_in_bits(PE_11_io_data_1_in_bits),
    .io_data_1_out_valid(PE_11_io_data_1_out_valid),
    .io_data_1_out_bits(PE_11_io_data_1_out_bits),
    .io_data_0_in_valid(PE_11_io_data_0_in_valid),
    .io_data_0_in_bits(PE_11_io_data_0_in_bits),
    .io_data_0_out_valid(PE_11_io_data_0_out_valid),
    .io_data_0_out_bits(PE_11_io_data_0_out_bits),
    .io_sig_stat2trans(PE_11_io_sig_stat2trans)
  );
  PE PE_12 ( // @[pearray.scala 101:13]
    .clock(PE_12_clock),
    .reset(PE_12_reset),
    .io_data_2_in_bits(PE_12_io_data_2_in_bits),
    .io_data_2_out_bits(PE_12_io_data_2_out_bits),
    .io_data_1_in_valid(PE_12_io_data_1_in_valid),
    .io_data_1_in_bits(PE_12_io_data_1_in_bits),
    .io_data_1_out_valid(PE_12_io_data_1_out_valid),
    .io_data_1_out_bits(PE_12_io_data_1_out_bits),
    .io_data_0_in_valid(PE_12_io_data_0_in_valid),
    .io_data_0_in_bits(PE_12_io_data_0_in_bits),
    .io_data_0_out_valid(PE_12_io_data_0_out_valid),
    .io_data_0_out_bits(PE_12_io_data_0_out_bits),
    .io_sig_stat2trans(PE_12_io_sig_stat2trans)
  );
  PE PE_13 ( // @[pearray.scala 101:13]
    .clock(PE_13_clock),
    .reset(PE_13_reset),
    .io_data_2_in_bits(PE_13_io_data_2_in_bits),
    .io_data_2_out_bits(PE_13_io_data_2_out_bits),
    .io_data_1_in_valid(PE_13_io_data_1_in_valid),
    .io_data_1_in_bits(PE_13_io_data_1_in_bits),
    .io_data_1_out_valid(PE_13_io_data_1_out_valid),
    .io_data_1_out_bits(PE_13_io_data_1_out_bits),
    .io_data_0_in_valid(PE_13_io_data_0_in_valid),
    .io_data_0_in_bits(PE_13_io_data_0_in_bits),
    .io_data_0_out_valid(PE_13_io_data_0_out_valid),
    .io_data_0_out_bits(PE_13_io_data_0_out_bits),
    .io_sig_stat2trans(PE_13_io_sig_stat2trans)
  );
  PE PE_14 ( // @[pearray.scala 101:13]
    .clock(PE_14_clock),
    .reset(PE_14_reset),
    .io_data_2_in_bits(PE_14_io_data_2_in_bits),
    .io_data_2_out_bits(PE_14_io_data_2_out_bits),
    .io_data_1_in_valid(PE_14_io_data_1_in_valid),
    .io_data_1_in_bits(PE_14_io_data_1_in_bits),
    .io_data_1_out_valid(PE_14_io_data_1_out_valid),
    .io_data_1_out_bits(PE_14_io_data_1_out_bits),
    .io_data_0_in_valid(PE_14_io_data_0_in_valid),
    .io_data_0_in_bits(PE_14_io_data_0_in_bits),
    .io_data_0_out_valid(PE_14_io_data_0_out_valid),
    .io_data_0_out_bits(PE_14_io_data_0_out_bits),
    .io_sig_stat2trans(PE_14_io_sig_stat2trans)
  );
  PE PE_15 ( // @[pearray.scala 101:13]
    .clock(PE_15_clock),
    .reset(PE_15_reset),
    .io_data_2_in_bits(PE_15_io_data_2_in_bits),
    .io_data_2_out_bits(PE_15_io_data_2_out_bits),
    .io_data_1_in_valid(PE_15_io_data_1_in_valid),
    .io_data_1_in_bits(PE_15_io_data_1_in_bits),
    .io_data_1_out_valid(PE_15_io_data_1_out_valid),
    .io_data_1_out_bits(PE_15_io_data_1_out_bits),
    .io_data_0_in_valid(PE_15_io_data_0_in_valid),
    .io_data_0_in_bits(PE_15_io_data_0_in_bits),
    .io_data_0_out_valid(PE_15_io_data_0_out_valid),
    .io_data_0_out_bits(PE_15_io_data_0_out_bits),
    .io_sig_stat2trans(PE_15_io_sig_stat2trans)
  );
  PE PE_16 ( // @[pearray.scala 101:13]
    .clock(PE_16_clock),
    .reset(PE_16_reset),
    .io_data_2_in_bits(PE_16_io_data_2_in_bits),
    .io_data_2_out_bits(PE_16_io_data_2_out_bits),
    .io_data_1_in_valid(PE_16_io_data_1_in_valid),
    .io_data_1_in_bits(PE_16_io_data_1_in_bits),
    .io_data_1_out_valid(PE_16_io_data_1_out_valid),
    .io_data_1_out_bits(PE_16_io_data_1_out_bits),
    .io_data_0_in_valid(PE_16_io_data_0_in_valid),
    .io_data_0_in_bits(PE_16_io_data_0_in_bits),
    .io_data_0_out_valid(PE_16_io_data_0_out_valid),
    .io_data_0_out_bits(PE_16_io_data_0_out_bits),
    .io_sig_stat2trans(PE_16_io_sig_stat2trans)
  );
  PE PE_17 ( // @[pearray.scala 101:13]
    .clock(PE_17_clock),
    .reset(PE_17_reset),
    .io_data_2_in_bits(PE_17_io_data_2_in_bits),
    .io_data_2_out_bits(PE_17_io_data_2_out_bits),
    .io_data_1_in_valid(PE_17_io_data_1_in_valid),
    .io_data_1_in_bits(PE_17_io_data_1_in_bits),
    .io_data_1_out_valid(PE_17_io_data_1_out_valid),
    .io_data_1_out_bits(PE_17_io_data_1_out_bits),
    .io_data_0_in_valid(PE_17_io_data_0_in_valid),
    .io_data_0_in_bits(PE_17_io_data_0_in_bits),
    .io_data_0_out_valid(PE_17_io_data_0_out_valid),
    .io_data_0_out_bits(PE_17_io_data_0_out_bits),
    .io_sig_stat2trans(PE_17_io_sig_stat2trans)
  );
  PE PE_18 ( // @[pearray.scala 101:13]
    .clock(PE_18_clock),
    .reset(PE_18_reset),
    .io_data_2_in_bits(PE_18_io_data_2_in_bits),
    .io_data_2_out_bits(PE_18_io_data_2_out_bits),
    .io_data_1_in_valid(PE_18_io_data_1_in_valid),
    .io_data_1_in_bits(PE_18_io_data_1_in_bits),
    .io_data_1_out_valid(PE_18_io_data_1_out_valid),
    .io_data_1_out_bits(PE_18_io_data_1_out_bits),
    .io_data_0_in_valid(PE_18_io_data_0_in_valid),
    .io_data_0_in_bits(PE_18_io_data_0_in_bits),
    .io_data_0_out_valid(PE_18_io_data_0_out_valid),
    .io_data_0_out_bits(PE_18_io_data_0_out_bits),
    .io_sig_stat2trans(PE_18_io_sig_stat2trans)
  );
  PE PE_19 ( // @[pearray.scala 101:13]
    .clock(PE_19_clock),
    .reset(PE_19_reset),
    .io_data_2_in_bits(PE_19_io_data_2_in_bits),
    .io_data_2_out_bits(PE_19_io_data_2_out_bits),
    .io_data_1_in_valid(PE_19_io_data_1_in_valid),
    .io_data_1_in_bits(PE_19_io_data_1_in_bits),
    .io_data_1_out_valid(PE_19_io_data_1_out_valid),
    .io_data_1_out_bits(PE_19_io_data_1_out_bits),
    .io_data_0_in_valid(PE_19_io_data_0_in_valid),
    .io_data_0_in_bits(PE_19_io_data_0_in_bits),
    .io_data_0_out_valid(PE_19_io_data_0_out_valid),
    .io_data_0_out_bits(PE_19_io_data_0_out_bits),
    .io_sig_stat2trans(PE_19_io_sig_stat2trans)
  );
  PE PE_20 ( // @[pearray.scala 101:13]
    .clock(PE_20_clock),
    .reset(PE_20_reset),
    .io_data_2_in_bits(PE_20_io_data_2_in_bits),
    .io_data_2_out_bits(PE_20_io_data_2_out_bits),
    .io_data_1_in_valid(PE_20_io_data_1_in_valid),
    .io_data_1_in_bits(PE_20_io_data_1_in_bits),
    .io_data_1_out_valid(PE_20_io_data_1_out_valid),
    .io_data_1_out_bits(PE_20_io_data_1_out_bits),
    .io_data_0_in_valid(PE_20_io_data_0_in_valid),
    .io_data_0_in_bits(PE_20_io_data_0_in_bits),
    .io_data_0_out_valid(PE_20_io_data_0_out_valid),
    .io_data_0_out_bits(PE_20_io_data_0_out_bits),
    .io_sig_stat2trans(PE_20_io_sig_stat2trans)
  );
  PE PE_21 ( // @[pearray.scala 101:13]
    .clock(PE_21_clock),
    .reset(PE_21_reset),
    .io_data_2_in_bits(PE_21_io_data_2_in_bits),
    .io_data_2_out_bits(PE_21_io_data_2_out_bits),
    .io_data_1_in_valid(PE_21_io_data_1_in_valid),
    .io_data_1_in_bits(PE_21_io_data_1_in_bits),
    .io_data_1_out_valid(PE_21_io_data_1_out_valid),
    .io_data_1_out_bits(PE_21_io_data_1_out_bits),
    .io_data_0_in_valid(PE_21_io_data_0_in_valid),
    .io_data_0_in_bits(PE_21_io_data_0_in_bits),
    .io_data_0_out_valid(PE_21_io_data_0_out_valid),
    .io_data_0_out_bits(PE_21_io_data_0_out_bits),
    .io_sig_stat2trans(PE_21_io_sig_stat2trans)
  );
  PE PE_22 ( // @[pearray.scala 101:13]
    .clock(PE_22_clock),
    .reset(PE_22_reset),
    .io_data_2_in_bits(PE_22_io_data_2_in_bits),
    .io_data_2_out_bits(PE_22_io_data_2_out_bits),
    .io_data_1_in_valid(PE_22_io_data_1_in_valid),
    .io_data_1_in_bits(PE_22_io_data_1_in_bits),
    .io_data_1_out_valid(PE_22_io_data_1_out_valid),
    .io_data_1_out_bits(PE_22_io_data_1_out_bits),
    .io_data_0_in_valid(PE_22_io_data_0_in_valid),
    .io_data_0_in_bits(PE_22_io_data_0_in_bits),
    .io_data_0_out_valid(PE_22_io_data_0_out_valid),
    .io_data_0_out_bits(PE_22_io_data_0_out_bits),
    .io_sig_stat2trans(PE_22_io_sig_stat2trans)
  );
  PE PE_23 ( // @[pearray.scala 101:13]
    .clock(PE_23_clock),
    .reset(PE_23_reset),
    .io_data_2_in_bits(PE_23_io_data_2_in_bits),
    .io_data_2_out_bits(PE_23_io_data_2_out_bits),
    .io_data_1_in_valid(PE_23_io_data_1_in_valid),
    .io_data_1_in_bits(PE_23_io_data_1_in_bits),
    .io_data_1_out_valid(PE_23_io_data_1_out_valid),
    .io_data_1_out_bits(PE_23_io_data_1_out_bits),
    .io_data_0_in_valid(PE_23_io_data_0_in_valid),
    .io_data_0_in_bits(PE_23_io_data_0_in_bits),
    .io_data_0_out_valid(PE_23_io_data_0_out_valid),
    .io_data_0_out_bits(PE_23_io_data_0_out_bits),
    .io_sig_stat2trans(PE_23_io_sig_stat2trans)
  );
  PE PE_24 ( // @[pearray.scala 101:13]
    .clock(PE_24_clock),
    .reset(PE_24_reset),
    .io_data_2_in_bits(PE_24_io_data_2_in_bits),
    .io_data_2_out_bits(PE_24_io_data_2_out_bits),
    .io_data_1_in_valid(PE_24_io_data_1_in_valid),
    .io_data_1_in_bits(PE_24_io_data_1_in_bits),
    .io_data_1_out_valid(PE_24_io_data_1_out_valid),
    .io_data_1_out_bits(PE_24_io_data_1_out_bits),
    .io_data_0_in_valid(PE_24_io_data_0_in_valid),
    .io_data_0_in_bits(PE_24_io_data_0_in_bits),
    .io_data_0_out_valid(PE_24_io_data_0_out_valid),
    .io_data_0_out_bits(PE_24_io_data_0_out_bits),
    .io_sig_stat2trans(PE_24_io_sig_stat2trans)
  );
  PE PE_25 ( // @[pearray.scala 101:13]
    .clock(PE_25_clock),
    .reset(PE_25_reset),
    .io_data_2_in_bits(PE_25_io_data_2_in_bits),
    .io_data_2_out_bits(PE_25_io_data_2_out_bits),
    .io_data_1_in_valid(PE_25_io_data_1_in_valid),
    .io_data_1_in_bits(PE_25_io_data_1_in_bits),
    .io_data_1_out_valid(PE_25_io_data_1_out_valid),
    .io_data_1_out_bits(PE_25_io_data_1_out_bits),
    .io_data_0_in_valid(PE_25_io_data_0_in_valid),
    .io_data_0_in_bits(PE_25_io_data_0_in_bits),
    .io_data_0_out_valid(PE_25_io_data_0_out_valid),
    .io_data_0_out_bits(PE_25_io_data_0_out_bits),
    .io_sig_stat2trans(PE_25_io_sig_stat2trans)
  );
  PE PE_26 ( // @[pearray.scala 101:13]
    .clock(PE_26_clock),
    .reset(PE_26_reset),
    .io_data_2_in_bits(PE_26_io_data_2_in_bits),
    .io_data_2_out_bits(PE_26_io_data_2_out_bits),
    .io_data_1_in_valid(PE_26_io_data_1_in_valid),
    .io_data_1_in_bits(PE_26_io_data_1_in_bits),
    .io_data_1_out_valid(PE_26_io_data_1_out_valid),
    .io_data_1_out_bits(PE_26_io_data_1_out_bits),
    .io_data_0_in_valid(PE_26_io_data_0_in_valid),
    .io_data_0_in_bits(PE_26_io_data_0_in_bits),
    .io_data_0_out_valid(PE_26_io_data_0_out_valid),
    .io_data_0_out_bits(PE_26_io_data_0_out_bits),
    .io_sig_stat2trans(PE_26_io_sig_stat2trans)
  );
  PE PE_27 ( // @[pearray.scala 101:13]
    .clock(PE_27_clock),
    .reset(PE_27_reset),
    .io_data_2_in_bits(PE_27_io_data_2_in_bits),
    .io_data_2_out_bits(PE_27_io_data_2_out_bits),
    .io_data_1_in_valid(PE_27_io_data_1_in_valid),
    .io_data_1_in_bits(PE_27_io_data_1_in_bits),
    .io_data_1_out_valid(PE_27_io_data_1_out_valid),
    .io_data_1_out_bits(PE_27_io_data_1_out_bits),
    .io_data_0_in_valid(PE_27_io_data_0_in_valid),
    .io_data_0_in_bits(PE_27_io_data_0_in_bits),
    .io_data_0_out_valid(PE_27_io_data_0_out_valid),
    .io_data_0_out_bits(PE_27_io_data_0_out_bits),
    .io_sig_stat2trans(PE_27_io_sig_stat2trans)
  );
  PE PE_28 ( // @[pearray.scala 101:13]
    .clock(PE_28_clock),
    .reset(PE_28_reset),
    .io_data_2_in_bits(PE_28_io_data_2_in_bits),
    .io_data_2_out_bits(PE_28_io_data_2_out_bits),
    .io_data_1_in_valid(PE_28_io_data_1_in_valid),
    .io_data_1_in_bits(PE_28_io_data_1_in_bits),
    .io_data_1_out_valid(PE_28_io_data_1_out_valid),
    .io_data_1_out_bits(PE_28_io_data_1_out_bits),
    .io_data_0_in_valid(PE_28_io_data_0_in_valid),
    .io_data_0_in_bits(PE_28_io_data_0_in_bits),
    .io_data_0_out_valid(PE_28_io_data_0_out_valid),
    .io_data_0_out_bits(PE_28_io_data_0_out_bits),
    .io_sig_stat2trans(PE_28_io_sig_stat2trans)
  );
  PE PE_29 ( // @[pearray.scala 101:13]
    .clock(PE_29_clock),
    .reset(PE_29_reset),
    .io_data_2_in_bits(PE_29_io_data_2_in_bits),
    .io_data_2_out_bits(PE_29_io_data_2_out_bits),
    .io_data_1_in_valid(PE_29_io_data_1_in_valid),
    .io_data_1_in_bits(PE_29_io_data_1_in_bits),
    .io_data_1_out_valid(PE_29_io_data_1_out_valid),
    .io_data_1_out_bits(PE_29_io_data_1_out_bits),
    .io_data_0_in_valid(PE_29_io_data_0_in_valid),
    .io_data_0_in_bits(PE_29_io_data_0_in_bits),
    .io_data_0_out_valid(PE_29_io_data_0_out_valid),
    .io_data_0_out_bits(PE_29_io_data_0_out_bits),
    .io_sig_stat2trans(PE_29_io_sig_stat2trans)
  );
  PE PE_30 ( // @[pearray.scala 101:13]
    .clock(PE_30_clock),
    .reset(PE_30_reset),
    .io_data_2_in_bits(PE_30_io_data_2_in_bits),
    .io_data_2_out_bits(PE_30_io_data_2_out_bits),
    .io_data_1_in_valid(PE_30_io_data_1_in_valid),
    .io_data_1_in_bits(PE_30_io_data_1_in_bits),
    .io_data_1_out_valid(PE_30_io_data_1_out_valid),
    .io_data_1_out_bits(PE_30_io_data_1_out_bits),
    .io_data_0_in_valid(PE_30_io_data_0_in_valid),
    .io_data_0_in_bits(PE_30_io_data_0_in_bits),
    .io_data_0_out_valid(PE_30_io_data_0_out_valid),
    .io_data_0_out_bits(PE_30_io_data_0_out_bits),
    .io_sig_stat2trans(PE_30_io_sig_stat2trans)
  );
  PE PE_31 ( // @[pearray.scala 101:13]
    .clock(PE_31_clock),
    .reset(PE_31_reset),
    .io_data_2_in_bits(PE_31_io_data_2_in_bits),
    .io_data_2_out_bits(PE_31_io_data_2_out_bits),
    .io_data_1_in_valid(PE_31_io_data_1_in_valid),
    .io_data_1_in_bits(PE_31_io_data_1_in_bits),
    .io_data_1_out_valid(PE_31_io_data_1_out_valid),
    .io_data_1_out_bits(PE_31_io_data_1_out_bits),
    .io_data_0_in_valid(PE_31_io_data_0_in_valid),
    .io_data_0_in_bits(PE_31_io_data_0_in_bits),
    .io_data_0_out_valid(PE_31_io_data_0_out_valid),
    .io_data_0_out_bits(PE_31_io_data_0_out_bits),
    .io_sig_stat2trans(PE_31_io_sig_stat2trans)
  );
  PE PE_32 ( // @[pearray.scala 101:13]
    .clock(PE_32_clock),
    .reset(PE_32_reset),
    .io_data_2_in_bits(PE_32_io_data_2_in_bits),
    .io_data_2_out_bits(PE_32_io_data_2_out_bits),
    .io_data_1_in_valid(PE_32_io_data_1_in_valid),
    .io_data_1_in_bits(PE_32_io_data_1_in_bits),
    .io_data_1_out_valid(PE_32_io_data_1_out_valid),
    .io_data_1_out_bits(PE_32_io_data_1_out_bits),
    .io_data_0_in_valid(PE_32_io_data_0_in_valid),
    .io_data_0_in_bits(PE_32_io_data_0_in_bits),
    .io_data_0_out_valid(PE_32_io_data_0_out_valid),
    .io_data_0_out_bits(PE_32_io_data_0_out_bits),
    .io_sig_stat2trans(PE_32_io_sig_stat2trans)
  );
  PE PE_33 ( // @[pearray.scala 101:13]
    .clock(PE_33_clock),
    .reset(PE_33_reset),
    .io_data_2_in_bits(PE_33_io_data_2_in_bits),
    .io_data_2_out_bits(PE_33_io_data_2_out_bits),
    .io_data_1_in_valid(PE_33_io_data_1_in_valid),
    .io_data_1_in_bits(PE_33_io_data_1_in_bits),
    .io_data_1_out_valid(PE_33_io_data_1_out_valid),
    .io_data_1_out_bits(PE_33_io_data_1_out_bits),
    .io_data_0_in_valid(PE_33_io_data_0_in_valid),
    .io_data_0_in_bits(PE_33_io_data_0_in_bits),
    .io_data_0_out_valid(PE_33_io_data_0_out_valid),
    .io_data_0_out_bits(PE_33_io_data_0_out_bits),
    .io_sig_stat2trans(PE_33_io_sig_stat2trans)
  );
  PE PE_34 ( // @[pearray.scala 101:13]
    .clock(PE_34_clock),
    .reset(PE_34_reset),
    .io_data_2_in_bits(PE_34_io_data_2_in_bits),
    .io_data_2_out_bits(PE_34_io_data_2_out_bits),
    .io_data_1_in_valid(PE_34_io_data_1_in_valid),
    .io_data_1_in_bits(PE_34_io_data_1_in_bits),
    .io_data_1_out_valid(PE_34_io_data_1_out_valid),
    .io_data_1_out_bits(PE_34_io_data_1_out_bits),
    .io_data_0_in_valid(PE_34_io_data_0_in_valid),
    .io_data_0_in_bits(PE_34_io_data_0_in_bits),
    .io_data_0_out_valid(PE_34_io_data_0_out_valid),
    .io_data_0_out_bits(PE_34_io_data_0_out_bits),
    .io_sig_stat2trans(PE_34_io_sig_stat2trans)
  );
  PE PE_35 ( // @[pearray.scala 101:13]
    .clock(PE_35_clock),
    .reset(PE_35_reset),
    .io_data_2_in_bits(PE_35_io_data_2_in_bits),
    .io_data_2_out_bits(PE_35_io_data_2_out_bits),
    .io_data_1_in_valid(PE_35_io_data_1_in_valid),
    .io_data_1_in_bits(PE_35_io_data_1_in_bits),
    .io_data_1_out_valid(PE_35_io_data_1_out_valid),
    .io_data_1_out_bits(PE_35_io_data_1_out_bits),
    .io_data_0_in_valid(PE_35_io_data_0_in_valid),
    .io_data_0_in_bits(PE_35_io_data_0_in_bits),
    .io_data_0_out_valid(PE_35_io_data_0_out_valid),
    .io_data_0_out_bits(PE_35_io_data_0_out_bits),
    .io_sig_stat2trans(PE_35_io_sig_stat2trans)
  );
  PE PE_36 ( // @[pearray.scala 101:13]
    .clock(PE_36_clock),
    .reset(PE_36_reset),
    .io_data_2_in_bits(PE_36_io_data_2_in_bits),
    .io_data_2_out_bits(PE_36_io_data_2_out_bits),
    .io_data_1_in_valid(PE_36_io_data_1_in_valid),
    .io_data_1_in_bits(PE_36_io_data_1_in_bits),
    .io_data_1_out_valid(PE_36_io_data_1_out_valid),
    .io_data_1_out_bits(PE_36_io_data_1_out_bits),
    .io_data_0_in_valid(PE_36_io_data_0_in_valid),
    .io_data_0_in_bits(PE_36_io_data_0_in_bits),
    .io_data_0_out_valid(PE_36_io_data_0_out_valid),
    .io_data_0_out_bits(PE_36_io_data_0_out_bits),
    .io_sig_stat2trans(PE_36_io_sig_stat2trans)
  );
  PE PE_37 ( // @[pearray.scala 101:13]
    .clock(PE_37_clock),
    .reset(PE_37_reset),
    .io_data_2_in_bits(PE_37_io_data_2_in_bits),
    .io_data_2_out_bits(PE_37_io_data_2_out_bits),
    .io_data_1_in_valid(PE_37_io_data_1_in_valid),
    .io_data_1_in_bits(PE_37_io_data_1_in_bits),
    .io_data_1_out_valid(PE_37_io_data_1_out_valid),
    .io_data_1_out_bits(PE_37_io_data_1_out_bits),
    .io_data_0_in_valid(PE_37_io_data_0_in_valid),
    .io_data_0_in_bits(PE_37_io_data_0_in_bits),
    .io_data_0_out_valid(PE_37_io_data_0_out_valid),
    .io_data_0_out_bits(PE_37_io_data_0_out_bits),
    .io_sig_stat2trans(PE_37_io_sig_stat2trans)
  );
  PE PE_38 ( // @[pearray.scala 101:13]
    .clock(PE_38_clock),
    .reset(PE_38_reset),
    .io_data_2_in_bits(PE_38_io_data_2_in_bits),
    .io_data_2_out_bits(PE_38_io_data_2_out_bits),
    .io_data_1_in_valid(PE_38_io_data_1_in_valid),
    .io_data_1_in_bits(PE_38_io_data_1_in_bits),
    .io_data_1_out_valid(PE_38_io_data_1_out_valid),
    .io_data_1_out_bits(PE_38_io_data_1_out_bits),
    .io_data_0_in_valid(PE_38_io_data_0_in_valid),
    .io_data_0_in_bits(PE_38_io_data_0_in_bits),
    .io_data_0_out_valid(PE_38_io_data_0_out_valid),
    .io_data_0_out_bits(PE_38_io_data_0_out_bits),
    .io_sig_stat2trans(PE_38_io_sig_stat2trans)
  );
  PE PE_39 ( // @[pearray.scala 101:13]
    .clock(PE_39_clock),
    .reset(PE_39_reset),
    .io_data_2_in_bits(PE_39_io_data_2_in_bits),
    .io_data_2_out_bits(PE_39_io_data_2_out_bits),
    .io_data_1_in_valid(PE_39_io_data_1_in_valid),
    .io_data_1_in_bits(PE_39_io_data_1_in_bits),
    .io_data_1_out_valid(PE_39_io_data_1_out_valid),
    .io_data_1_out_bits(PE_39_io_data_1_out_bits),
    .io_data_0_in_valid(PE_39_io_data_0_in_valid),
    .io_data_0_in_bits(PE_39_io_data_0_in_bits),
    .io_data_0_out_valid(PE_39_io_data_0_out_valid),
    .io_data_0_out_bits(PE_39_io_data_0_out_bits),
    .io_sig_stat2trans(PE_39_io_sig_stat2trans)
  );
  PE PE_40 ( // @[pearray.scala 101:13]
    .clock(PE_40_clock),
    .reset(PE_40_reset),
    .io_data_2_in_bits(PE_40_io_data_2_in_bits),
    .io_data_2_out_bits(PE_40_io_data_2_out_bits),
    .io_data_1_in_valid(PE_40_io_data_1_in_valid),
    .io_data_1_in_bits(PE_40_io_data_1_in_bits),
    .io_data_1_out_valid(PE_40_io_data_1_out_valid),
    .io_data_1_out_bits(PE_40_io_data_1_out_bits),
    .io_data_0_in_valid(PE_40_io_data_0_in_valid),
    .io_data_0_in_bits(PE_40_io_data_0_in_bits),
    .io_data_0_out_valid(PE_40_io_data_0_out_valid),
    .io_data_0_out_bits(PE_40_io_data_0_out_bits),
    .io_sig_stat2trans(PE_40_io_sig_stat2trans)
  );
  PE PE_41 ( // @[pearray.scala 101:13]
    .clock(PE_41_clock),
    .reset(PE_41_reset),
    .io_data_2_in_bits(PE_41_io_data_2_in_bits),
    .io_data_2_out_bits(PE_41_io_data_2_out_bits),
    .io_data_1_in_valid(PE_41_io_data_1_in_valid),
    .io_data_1_in_bits(PE_41_io_data_1_in_bits),
    .io_data_1_out_valid(PE_41_io_data_1_out_valid),
    .io_data_1_out_bits(PE_41_io_data_1_out_bits),
    .io_data_0_in_valid(PE_41_io_data_0_in_valid),
    .io_data_0_in_bits(PE_41_io_data_0_in_bits),
    .io_data_0_out_valid(PE_41_io_data_0_out_valid),
    .io_data_0_out_bits(PE_41_io_data_0_out_bits),
    .io_sig_stat2trans(PE_41_io_sig_stat2trans)
  );
  PE PE_42 ( // @[pearray.scala 101:13]
    .clock(PE_42_clock),
    .reset(PE_42_reset),
    .io_data_2_in_bits(PE_42_io_data_2_in_bits),
    .io_data_2_out_bits(PE_42_io_data_2_out_bits),
    .io_data_1_in_valid(PE_42_io_data_1_in_valid),
    .io_data_1_in_bits(PE_42_io_data_1_in_bits),
    .io_data_1_out_valid(PE_42_io_data_1_out_valid),
    .io_data_1_out_bits(PE_42_io_data_1_out_bits),
    .io_data_0_in_valid(PE_42_io_data_0_in_valid),
    .io_data_0_in_bits(PE_42_io_data_0_in_bits),
    .io_data_0_out_valid(PE_42_io_data_0_out_valid),
    .io_data_0_out_bits(PE_42_io_data_0_out_bits),
    .io_sig_stat2trans(PE_42_io_sig_stat2trans)
  );
  PE PE_43 ( // @[pearray.scala 101:13]
    .clock(PE_43_clock),
    .reset(PE_43_reset),
    .io_data_2_in_bits(PE_43_io_data_2_in_bits),
    .io_data_2_out_bits(PE_43_io_data_2_out_bits),
    .io_data_1_in_valid(PE_43_io_data_1_in_valid),
    .io_data_1_in_bits(PE_43_io_data_1_in_bits),
    .io_data_1_out_valid(PE_43_io_data_1_out_valid),
    .io_data_1_out_bits(PE_43_io_data_1_out_bits),
    .io_data_0_in_valid(PE_43_io_data_0_in_valid),
    .io_data_0_in_bits(PE_43_io_data_0_in_bits),
    .io_data_0_out_valid(PE_43_io_data_0_out_valid),
    .io_data_0_out_bits(PE_43_io_data_0_out_bits),
    .io_sig_stat2trans(PE_43_io_sig_stat2trans)
  );
  PE PE_44 ( // @[pearray.scala 101:13]
    .clock(PE_44_clock),
    .reset(PE_44_reset),
    .io_data_2_in_bits(PE_44_io_data_2_in_bits),
    .io_data_2_out_bits(PE_44_io_data_2_out_bits),
    .io_data_1_in_valid(PE_44_io_data_1_in_valid),
    .io_data_1_in_bits(PE_44_io_data_1_in_bits),
    .io_data_1_out_valid(PE_44_io_data_1_out_valid),
    .io_data_1_out_bits(PE_44_io_data_1_out_bits),
    .io_data_0_in_valid(PE_44_io_data_0_in_valid),
    .io_data_0_in_bits(PE_44_io_data_0_in_bits),
    .io_data_0_out_valid(PE_44_io_data_0_out_valid),
    .io_data_0_out_bits(PE_44_io_data_0_out_bits),
    .io_sig_stat2trans(PE_44_io_sig_stat2trans)
  );
  PE PE_45 ( // @[pearray.scala 101:13]
    .clock(PE_45_clock),
    .reset(PE_45_reset),
    .io_data_2_in_bits(PE_45_io_data_2_in_bits),
    .io_data_2_out_bits(PE_45_io_data_2_out_bits),
    .io_data_1_in_valid(PE_45_io_data_1_in_valid),
    .io_data_1_in_bits(PE_45_io_data_1_in_bits),
    .io_data_1_out_valid(PE_45_io_data_1_out_valid),
    .io_data_1_out_bits(PE_45_io_data_1_out_bits),
    .io_data_0_in_valid(PE_45_io_data_0_in_valid),
    .io_data_0_in_bits(PE_45_io_data_0_in_bits),
    .io_data_0_out_valid(PE_45_io_data_0_out_valid),
    .io_data_0_out_bits(PE_45_io_data_0_out_bits),
    .io_sig_stat2trans(PE_45_io_sig_stat2trans)
  );
  PE PE_46 ( // @[pearray.scala 101:13]
    .clock(PE_46_clock),
    .reset(PE_46_reset),
    .io_data_2_in_bits(PE_46_io_data_2_in_bits),
    .io_data_2_out_bits(PE_46_io_data_2_out_bits),
    .io_data_1_in_valid(PE_46_io_data_1_in_valid),
    .io_data_1_in_bits(PE_46_io_data_1_in_bits),
    .io_data_1_out_valid(PE_46_io_data_1_out_valid),
    .io_data_1_out_bits(PE_46_io_data_1_out_bits),
    .io_data_0_in_valid(PE_46_io_data_0_in_valid),
    .io_data_0_in_bits(PE_46_io_data_0_in_bits),
    .io_data_0_out_valid(PE_46_io_data_0_out_valid),
    .io_data_0_out_bits(PE_46_io_data_0_out_bits),
    .io_sig_stat2trans(PE_46_io_sig_stat2trans)
  );
  PE PE_47 ( // @[pearray.scala 101:13]
    .clock(PE_47_clock),
    .reset(PE_47_reset),
    .io_data_2_in_bits(PE_47_io_data_2_in_bits),
    .io_data_2_out_bits(PE_47_io_data_2_out_bits),
    .io_data_1_in_valid(PE_47_io_data_1_in_valid),
    .io_data_1_in_bits(PE_47_io_data_1_in_bits),
    .io_data_1_out_valid(PE_47_io_data_1_out_valid),
    .io_data_1_out_bits(PE_47_io_data_1_out_bits),
    .io_data_0_in_valid(PE_47_io_data_0_in_valid),
    .io_data_0_in_bits(PE_47_io_data_0_in_bits),
    .io_data_0_out_valid(PE_47_io_data_0_out_valid),
    .io_data_0_out_bits(PE_47_io_data_0_out_bits),
    .io_sig_stat2trans(PE_47_io_sig_stat2trans)
  );
  PE PE_48 ( // @[pearray.scala 101:13]
    .clock(PE_48_clock),
    .reset(PE_48_reset),
    .io_data_2_in_bits(PE_48_io_data_2_in_bits),
    .io_data_2_out_bits(PE_48_io_data_2_out_bits),
    .io_data_1_in_valid(PE_48_io_data_1_in_valid),
    .io_data_1_in_bits(PE_48_io_data_1_in_bits),
    .io_data_1_out_valid(PE_48_io_data_1_out_valid),
    .io_data_1_out_bits(PE_48_io_data_1_out_bits),
    .io_data_0_in_valid(PE_48_io_data_0_in_valid),
    .io_data_0_in_bits(PE_48_io_data_0_in_bits),
    .io_data_0_out_valid(PE_48_io_data_0_out_valid),
    .io_data_0_out_bits(PE_48_io_data_0_out_bits),
    .io_sig_stat2trans(PE_48_io_sig_stat2trans)
  );
  PE PE_49 ( // @[pearray.scala 101:13]
    .clock(PE_49_clock),
    .reset(PE_49_reset),
    .io_data_2_in_bits(PE_49_io_data_2_in_bits),
    .io_data_2_out_bits(PE_49_io_data_2_out_bits),
    .io_data_1_in_valid(PE_49_io_data_1_in_valid),
    .io_data_1_in_bits(PE_49_io_data_1_in_bits),
    .io_data_1_out_valid(PE_49_io_data_1_out_valid),
    .io_data_1_out_bits(PE_49_io_data_1_out_bits),
    .io_data_0_in_valid(PE_49_io_data_0_in_valid),
    .io_data_0_in_bits(PE_49_io_data_0_in_bits),
    .io_data_0_out_valid(PE_49_io_data_0_out_valid),
    .io_data_0_out_bits(PE_49_io_data_0_out_bits),
    .io_sig_stat2trans(PE_49_io_sig_stat2trans)
  );
  PE PE_50 ( // @[pearray.scala 101:13]
    .clock(PE_50_clock),
    .reset(PE_50_reset),
    .io_data_2_in_bits(PE_50_io_data_2_in_bits),
    .io_data_2_out_bits(PE_50_io_data_2_out_bits),
    .io_data_1_in_valid(PE_50_io_data_1_in_valid),
    .io_data_1_in_bits(PE_50_io_data_1_in_bits),
    .io_data_1_out_valid(PE_50_io_data_1_out_valid),
    .io_data_1_out_bits(PE_50_io_data_1_out_bits),
    .io_data_0_in_valid(PE_50_io_data_0_in_valid),
    .io_data_0_in_bits(PE_50_io_data_0_in_bits),
    .io_data_0_out_valid(PE_50_io_data_0_out_valid),
    .io_data_0_out_bits(PE_50_io_data_0_out_bits),
    .io_sig_stat2trans(PE_50_io_sig_stat2trans)
  );
  PE PE_51 ( // @[pearray.scala 101:13]
    .clock(PE_51_clock),
    .reset(PE_51_reset),
    .io_data_2_in_bits(PE_51_io_data_2_in_bits),
    .io_data_2_out_bits(PE_51_io_data_2_out_bits),
    .io_data_1_in_valid(PE_51_io_data_1_in_valid),
    .io_data_1_in_bits(PE_51_io_data_1_in_bits),
    .io_data_1_out_valid(PE_51_io_data_1_out_valid),
    .io_data_1_out_bits(PE_51_io_data_1_out_bits),
    .io_data_0_in_valid(PE_51_io_data_0_in_valid),
    .io_data_0_in_bits(PE_51_io_data_0_in_bits),
    .io_data_0_out_valid(PE_51_io_data_0_out_valid),
    .io_data_0_out_bits(PE_51_io_data_0_out_bits),
    .io_sig_stat2trans(PE_51_io_sig_stat2trans)
  );
  PE PE_52 ( // @[pearray.scala 101:13]
    .clock(PE_52_clock),
    .reset(PE_52_reset),
    .io_data_2_in_bits(PE_52_io_data_2_in_bits),
    .io_data_2_out_bits(PE_52_io_data_2_out_bits),
    .io_data_1_in_valid(PE_52_io_data_1_in_valid),
    .io_data_1_in_bits(PE_52_io_data_1_in_bits),
    .io_data_1_out_valid(PE_52_io_data_1_out_valid),
    .io_data_1_out_bits(PE_52_io_data_1_out_bits),
    .io_data_0_in_valid(PE_52_io_data_0_in_valid),
    .io_data_0_in_bits(PE_52_io_data_0_in_bits),
    .io_data_0_out_valid(PE_52_io_data_0_out_valid),
    .io_data_0_out_bits(PE_52_io_data_0_out_bits),
    .io_sig_stat2trans(PE_52_io_sig_stat2trans)
  );
  PE PE_53 ( // @[pearray.scala 101:13]
    .clock(PE_53_clock),
    .reset(PE_53_reset),
    .io_data_2_in_bits(PE_53_io_data_2_in_bits),
    .io_data_2_out_bits(PE_53_io_data_2_out_bits),
    .io_data_1_in_valid(PE_53_io_data_1_in_valid),
    .io_data_1_in_bits(PE_53_io_data_1_in_bits),
    .io_data_1_out_valid(PE_53_io_data_1_out_valid),
    .io_data_1_out_bits(PE_53_io_data_1_out_bits),
    .io_data_0_in_valid(PE_53_io_data_0_in_valid),
    .io_data_0_in_bits(PE_53_io_data_0_in_bits),
    .io_data_0_out_valid(PE_53_io_data_0_out_valid),
    .io_data_0_out_bits(PE_53_io_data_0_out_bits),
    .io_sig_stat2trans(PE_53_io_sig_stat2trans)
  );
  PE PE_54 ( // @[pearray.scala 101:13]
    .clock(PE_54_clock),
    .reset(PE_54_reset),
    .io_data_2_in_bits(PE_54_io_data_2_in_bits),
    .io_data_2_out_bits(PE_54_io_data_2_out_bits),
    .io_data_1_in_valid(PE_54_io_data_1_in_valid),
    .io_data_1_in_bits(PE_54_io_data_1_in_bits),
    .io_data_1_out_valid(PE_54_io_data_1_out_valid),
    .io_data_1_out_bits(PE_54_io_data_1_out_bits),
    .io_data_0_in_valid(PE_54_io_data_0_in_valid),
    .io_data_0_in_bits(PE_54_io_data_0_in_bits),
    .io_data_0_out_valid(PE_54_io_data_0_out_valid),
    .io_data_0_out_bits(PE_54_io_data_0_out_bits),
    .io_sig_stat2trans(PE_54_io_sig_stat2trans)
  );
  PE PE_55 ( // @[pearray.scala 101:13]
    .clock(PE_55_clock),
    .reset(PE_55_reset),
    .io_data_2_in_bits(PE_55_io_data_2_in_bits),
    .io_data_2_out_bits(PE_55_io_data_2_out_bits),
    .io_data_1_in_valid(PE_55_io_data_1_in_valid),
    .io_data_1_in_bits(PE_55_io_data_1_in_bits),
    .io_data_1_out_valid(PE_55_io_data_1_out_valid),
    .io_data_1_out_bits(PE_55_io_data_1_out_bits),
    .io_data_0_in_valid(PE_55_io_data_0_in_valid),
    .io_data_0_in_bits(PE_55_io_data_0_in_bits),
    .io_data_0_out_valid(PE_55_io_data_0_out_valid),
    .io_data_0_out_bits(PE_55_io_data_0_out_bits),
    .io_sig_stat2trans(PE_55_io_sig_stat2trans)
  );
  PE PE_56 ( // @[pearray.scala 101:13]
    .clock(PE_56_clock),
    .reset(PE_56_reset),
    .io_data_2_in_bits(PE_56_io_data_2_in_bits),
    .io_data_2_out_bits(PE_56_io_data_2_out_bits),
    .io_data_1_in_valid(PE_56_io_data_1_in_valid),
    .io_data_1_in_bits(PE_56_io_data_1_in_bits),
    .io_data_1_out_valid(PE_56_io_data_1_out_valid),
    .io_data_1_out_bits(PE_56_io_data_1_out_bits),
    .io_data_0_in_valid(PE_56_io_data_0_in_valid),
    .io_data_0_in_bits(PE_56_io_data_0_in_bits),
    .io_data_0_out_valid(PE_56_io_data_0_out_valid),
    .io_data_0_out_bits(PE_56_io_data_0_out_bits),
    .io_sig_stat2trans(PE_56_io_sig_stat2trans)
  );
  PE PE_57 ( // @[pearray.scala 101:13]
    .clock(PE_57_clock),
    .reset(PE_57_reset),
    .io_data_2_in_bits(PE_57_io_data_2_in_bits),
    .io_data_2_out_bits(PE_57_io_data_2_out_bits),
    .io_data_1_in_valid(PE_57_io_data_1_in_valid),
    .io_data_1_in_bits(PE_57_io_data_1_in_bits),
    .io_data_1_out_valid(PE_57_io_data_1_out_valid),
    .io_data_1_out_bits(PE_57_io_data_1_out_bits),
    .io_data_0_in_valid(PE_57_io_data_0_in_valid),
    .io_data_0_in_bits(PE_57_io_data_0_in_bits),
    .io_data_0_out_valid(PE_57_io_data_0_out_valid),
    .io_data_0_out_bits(PE_57_io_data_0_out_bits),
    .io_sig_stat2trans(PE_57_io_sig_stat2trans)
  );
  PE PE_58 ( // @[pearray.scala 101:13]
    .clock(PE_58_clock),
    .reset(PE_58_reset),
    .io_data_2_in_bits(PE_58_io_data_2_in_bits),
    .io_data_2_out_bits(PE_58_io_data_2_out_bits),
    .io_data_1_in_valid(PE_58_io_data_1_in_valid),
    .io_data_1_in_bits(PE_58_io_data_1_in_bits),
    .io_data_1_out_valid(PE_58_io_data_1_out_valid),
    .io_data_1_out_bits(PE_58_io_data_1_out_bits),
    .io_data_0_in_valid(PE_58_io_data_0_in_valid),
    .io_data_0_in_bits(PE_58_io_data_0_in_bits),
    .io_data_0_out_valid(PE_58_io_data_0_out_valid),
    .io_data_0_out_bits(PE_58_io_data_0_out_bits),
    .io_sig_stat2trans(PE_58_io_sig_stat2trans)
  );
  PE PE_59 ( // @[pearray.scala 101:13]
    .clock(PE_59_clock),
    .reset(PE_59_reset),
    .io_data_2_in_bits(PE_59_io_data_2_in_bits),
    .io_data_2_out_bits(PE_59_io_data_2_out_bits),
    .io_data_1_in_valid(PE_59_io_data_1_in_valid),
    .io_data_1_in_bits(PE_59_io_data_1_in_bits),
    .io_data_1_out_valid(PE_59_io_data_1_out_valid),
    .io_data_1_out_bits(PE_59_io_data_1_out_bits),
    .io_data_0_in_valid(PE_59_io_data_0_in_valid),
    .io_data_0_in_bits(PE_59_io_data_0_in_bits),
    .io_data_0_out_valid(PE_59_io_data_0_out_valid),
    .io_data_0_out_bits(PE_59_io_data_0_out_bits),
    .io_sig_stat2trans(PE_59_io_sig_stat2trans)
  );
  PE PE_60 ( // @[pearray.scala 101:13]
    .clock(PE_60_clock),
    .reset(PE_60_reset),
    .io_data_2_in_bits(PE_60_io_data_2_in_bits),
    .io_data_2_out_bits(PE_60_io_data_2_out_bits),
    .io_data_1_in_valid(PE_60_io_data_1_in_valid),
    .io_data_1_in_bits(PE_60_io_data_1_in_bits),
    .io_data_1_out_valid(PE_60_io_data_1_out_valid),
    .io_data_1_out_bits(PE_60_io_data_1_out_bits),
    .io_data_0_in_valid(PE_60_io_data_0_in_valid),
    .io_data_0_in_bits(PE_60_io_data_0_in_bits),
    .io_data_0_out_valid(PE_60_io_data_0_out_valid),
    .io_data_0_out_bits(PE_60_io_data_0_out_bits),
    .io_sig_stat2trans(PE_60_io_sig_stat2trans)
  );
  PE PE_61 ( // @[pearray.scala 101:13]
    .clock(PE_61_clock),
    .reset(PE_61_reset),
    .io_data_2_in_bits(PE_61_io_data_2_in_bits),
    .io_data_2_out_bits(PE_61_io_data_2_out_bits),
    .io_data_1_in_valid(PE_61_io_data_1_in_valid),
    .io_data_1_in_bits(PE_61_io_data_1_in_bits),
    .io_data_1_out_valid(PE_61_io_data_1_out_valid),
    .io_data_1_out_bits(PE_61_io_data_1_out_bits),
    .io_data_0_in_valid(PE_61_io_data_0_in_valid),
    .io_data_0_in_bits(PE_61_io_data_0_in_bits),
    .io_data_0_out_valid(PE_61_io_data_0_out_valid),
    .io_data_0_out_bits(PE_61_io_data_0_out_bits),
    .io_sig_stat2trans(PE_61_io_sig_stat2trans)
  );
  PE PE_62 ( // @[pearray.scala 101:13]
    .clock(PE_62_clock),
    .reset(PE_62_reset),
    .io_data_2_in_bits(PE_62_io_data_2_in_bits),
    .io_data_2_out_bits(PE_62_io_data_2_out_bits),
    .io_data_1_in_valid(PE_62_io_data_1_in_valid),
    .io_data_1_in_bits(PE_62_io_data_1_in_bits),
    .io_data_1_out_valid(PE_62_io_data_1_out_valid),
    .io_data_1_out_bits(PE_62_io_data_1_out_bits),
    .io_data_0_in_valid(PE_62_io_data_0_in_valid),
    .io_data_0_in_bits(PE_62_io_data_0_in_bits),
    .io_data_0_out_valid(PE_62_io_data_0_out_valid),
    .io_data_0_out_bits(PE_62_io_data_0_out_bits),
    .io_sig_stat2trans(PE_62_io_sig_stat2trans)
  );
  PE PE_63 ( // @[pearray.scala 101:13]
    .clock(PE_63_clock),
    .reset(PE_63_reset),
    .io_data_2_in_bits(PE_63_io_data_2_in_bits),
    .io_data_2_out_bits(PE_63_io_data_2_out_bits),
    .io_data_1_in_valid(PE_63_io_data_1_in_valid),
    .io_data_1_in_bits(PE_63_io_data_1_in_bits),
    .io_data_1_out_valid(PE_63_io_data_1_out_valid),
    .io_data_1_out_bits(PE_63_io_data_1_out_bits),
    .io_data_0_in_valid(PE_63_io_data_0_in_valid),
    .io_data_0_in_bits(PE_63_io_data_0_in_bits),
    .io_data_0_out_valid(PE_63_io_data_0_out_valid),
    .io_data_0_out_bits(PE_63_io_data_0_out_bits),
    .io_sig_stat2trans(PE_63_io_sig_stat2trans)
  );
  PE PE_64 ( // @[pearray.scala 101:13]
    .clock(PE_64_clock),
    .reset(PE_64_reset),
    .io_data_2_in_bits(PE_64_io_data_2_in_bits),
    .io_data_2_out_bits(PE_64_io_data_2_out_bits),
    .io_data_1_in_valid(PE_64_io_data_1_in_valid),
    .io_data_1_in_bits(PE_64_io_data_1_in_bits),
    .io_data_1_out_valid(PE_64_io_data_1_out_valid),
    .io_data_1_out_bits(PE_64_io_data_1_out_bits),
    .io_data_0_in_valid(PE_64_io_data_0_in_valid),
    .io_data_0_in_bits(PE_64_io_data_0_in_bits),
    .io_data_0_out_valid(PE_64_io_data_0_out_valid),
    .io_data_0_out_bits(PE_64_io_data_0_out_bits),
    .io_sig_stat2trans(PE_64_io_sig_stat2trans)
  );
  PE PE_65 ( // @[pearray.scala 101:13]
    .clock(PE_65_clock),
    .reset(PE_65_reset),
    .io_data_2_in_bits(PE_65_io_data_2_in_bits),
    .io_data_2_out_bits(PE_65_io_data_2_out_bits),
    .io_data_1_in_valid(PE_65_io_data_1_in_valid),
    .io_data_1_in_bits(PE_65_io_data_1_in_bits),
    .io_data_1_out_valid(PE_65_io_data_1_out_valid),
    .io_data_1_out_bits(PE_65_io_data_1_out_bits),
    .io_data_0_in_valid(PE_65_io_data_0_in_valid),
    .io_data_0_in_bits(PE_65_io_data_0_in_bits),
    .io_data_0_out_valid(PE_65_io_data_0_out_valid),
    .io_data_0_out_bits(PE_65_io_data_0_out_bits),
    .io_sig_stat2trans(PE_65_io_sig_stat2trans)
  );
  PE PE_66 ( // @[pearray.scala 101:13]
    .clock(PE_66_clock),
    .reset(PE_66_reset),
    .io_data_2_in_bits(PE_66_io_data_2_in_bits),
    .io_data_2_out_bits(PE_66_io_data_2_out_bits),
    .io_data_1_in_valid(PE_66_io_data_1_in_valid),
    .io_data_1_in_bits(PE_66_io_data_1_in_bits),
    .io_data_1_out_valid(PE_66_io_data_1_out_valid),
    .io_data_1_out_bits(PE_66_io_data_1_out_bits),
    .io_data_0_in_valid(PE_66_io_data_0_in_valid),
    .io_data_0_in_bits(PE_66_io_data_0_in_bits),
    .io_data_0_out_valid(PE_66_io_data_0_out_valid),
    .io_data_0_out_bits(PE_66_io_data_0_out_bits),
    .io_sig_stat2trans(PE_66_io_sig_stat2trans)
  );
  PE PE_67 ( // @[pearray.scala 101:13]
    .clock(PE_67_clock),
    .reset(PE_67_reset),
    .io_data_2_in_bits(PE_67_io_data_2_in_bits),
    .io_data_2_out_bits(PE_67_io_data_2_out_bits),
    .io_data_1_in_valid(PE_67_io_data_1_in_valid),
    .io_data_1_in_bits(PE_67_io_data_1_in_bits),
    .io_data_1_out_valid(PE_67_io_data_1_out_valid),
    .io_data_1_out_bits(PE_67_io_data_1_out_bits),
    .io_data_0_in_valid(PE_67_io_data_0_in_valid),
    .io_data_0_in_bits(PE_67_io_data_0_in_bits),
    .io_data_0_out_valid(PE_67_io_data_0_out_valid),
    .io_data_0_out_bits(PE_67_io_data_0_out_bits),
    .io_sig_stat2trans(PE_67_io_sig_stat2trans)
  );
  PE PE_68 ( // @[pearray.scala 101:13]
    .clock(PE_68_clock),
    .reset(PE_68_reset),
    .io_data_2_in_bits(PE_68_io_data_2_in_bits),
    .io_data_2_out_bits(PE_68_io_data_2_out_bits),
    .io_data_1_in_valid(PE_68_io_data_1_in_valid),
    .io_data_1_in_bits(PE_68_io_data_1_in_bits),
    .io_data_1_out_valid(PE_68_io_data_1_out_valid),
    .io_data_1_out_bits(PE_68_io_data_1_out_bits),
    .io_data_0_in_valid(PE_68_io_data_0_in_valid),
    .io_data_0_in_bits(PE_68_io_data_0_in_bits),
    .io_data_0_out_valid(PE_68_io_data_0_out_valid),
    .io_data_0_out_bits(PE_68_io_data_0_out_bits),
    .io_sig_stat2trans(PE_68_io_sig_stat2trans)
  );
  PE PE_69 ( // @[pearray.scala 101:13]
    .clock(PE_69_clock),
    .reset(PE_69_reset),
    .io_data_2_in_bits(PE_69_io_data_2_in_bits),
    .io_data_2_out_bits(PE_69_io_data_2_out_bits),
    .io_data_1_in_valid(PE_69_io_data_1_in_valid),
    .io_data_1_in_bits(PE_69_io_data_1_in_bits),
    .io_data_1_out_valid(PE_69_io_data_1_out_valid),
    .io_data_1_out_bits(PE_69_io_data_1_out_bits),
    .io_data_0_in_valid(PE_69_io_data_0_in_valid),
    .io_data_0_in_bits(PE_69_io_data_0_in_bits),
    .io_data_0_out_valid(PE_69_io_data_0_out_valid),
    .io_data_0_out_bits(PE_69_io_data_0_out_bits),
    .io_sig_stat2trans(PE_69_io_sig_stat2trans)
  );
  PE PE_70 ( // @[pearray.scala 101:13]
    .clock(PE_70_clock),
    .reset(PE_70_reset),
    .io_data_2_in_bits(PE_70_io_data_2_in_bits),
    .io_data_2_out_bits(PE_70_io_data_2_out_bits),
    .io_data_1_in_valid(PE_70_io_data_1_in_valid),
    .io_data_1_in_bits(PE_70_io_data_1_in_bits),
    .io_data_1_out_valid(PE_70_io_data_1_out_valid),
    .io_data_1_out_bits(PE_70_io_data_1_out_bits),
    .io_data_0_in_valid(PE_70_io_data_0_in_valid),
    .io_data_0_in_bits(PE_70_io_data_0_in_bits),
    .io_data_0_out_valid(PE_70_io_data_0_out_valid),
    .io_data_0_out_bits(PE_70_io_data_0_out_bits),
    .io_sig_stat2trans(PE_70_io_sig_stat2trans)
  );
  PE PE_71 ( // @[pearray.scala 101:13]
    .clock(PE_71_clock),
    .reset(PE_71_reset),
    .io_data_2_in_bits(PE_71_io_data_2_in_bits),
    .io_data_2_out_bits(PE_71_io_data_2_out_bits),
    .io_data_1_in_valid(PE_71_io_data_1_in_valid),
    .io_data_1_in_bits(PE_71_io_data_1_in_bits),
    .io_data_1_out_valid(PE_71_io_data_1_out_valid),
    .io_data_1_out_bits(PE_71_io_data_1_out_bits),
    .io_data_0_in_valid(PE_71_io_data_0_in_valid),
    .io_data_0_in_bits(PE_71_io_data_0_in_bits),
    .io_data_0_out_valid(PE_71_io_data_0_out_valid),
    .io_data_0_out_bits(PE_71_io_data_0_out_bits),
    .io_sig_stat2trans(PE_71_io_sig_stat2trans)
  );
  PE PE_72 ( // @[pearray.scala 101:13]
    .clock(PE_72_clock),
    .reset(PE_72_reset),
    .io_data_2_in_bits(PE_72_io_data_2_in_bits),
    .io_data_2_out_bits(PE_72_io_data_2_out_bits),
    .io_data_1_in_valid(PE_72_io_data_1_in_valid),
    .io_data_1_in_bits(PE_72_io_data_1_in_bits),
    .io_data_1_out_valid(PE_72_io_data_1_out_valid),
    .io_data_1_out_bits(PE_72_io_data_1_out_bits),
    .io_data_0_in_valid(PE_72_io_data_0_in_valid),
    .io_data_0_in_bits(PE_72_io_data_0_in_bits),
    .io_data_0_out_valid(PE_72_io_data_0_out_valid),
    .io_data_0_out_bits(PE_72_io_data_0_out_bits),
    .io_sig_stat2trans(PE_72_io_sig_stat2trans)
  );
  PE PE_73 ( // @[pearray.scala 101:13]
    .clock(PE_73_clock),
    .reset(PE_73_reset),
    .io_data_2_in_bits(PE_73_io_data_2_in_bits),
    .io_data_2_out_bits(PE_73_io_data_2_out_bits),
    .io_data_1_in_valid(PE_73_io_data_1_in_valid),
    .io_data_1_in_bits(PE_73_io_data_1_in_bits),
    .io_data_1_out_valid(PE_73_io_data_1_out_valid),
    .io_data_1_out_bits(PE_73_io_data_1_out_bits),
    .io_data_0_in_valid(PE_73_io_data_0_in_valid),
    .io_data_0_in_bits(PE_73_io_data_0_in_bits),
    .io_data_0_out_valid(PE_73_io_data_0_out_valid),
    .io_data_0_out_bits(PE_73_io_data_0_out_bits),
    .io_sig_stat2trans(PE_73_io_sig_stat2trans)
  );
  PE PE_74 ( // @[pearray.scala 101:13]
    .clock(PE_74_clock),
    .reset(PE_74_reset),
    .io_data_2_in_bits(PE_74_io_data_2_in_bits),
    .io_data_2_out_bits(PE_74_io_data_2_out_bits),
    .io_data_1_in_valid(PE_74_io_data_1_in_valid),
    .io_data_1_in_bits(PE_74_io_data_1_in_bits),
    .io_data_1_out_valid(PE_74_io_data_1_out_valid),
    .io_data_1_out_bits(PE_74_io_data_1_out_bits),
    .io_data_0_in_valid(PE_74_io_data_0_in_valid),
    .io_data_0_in_bits(PE_74_io_data_0_in_bits),
    .io_data_0_out_valid(PE_74_io_data_0_out_valid),
    .io_data_0_out_bits(PE_74_io_data_0_out_bits),
    .io_sig_stat2trans(PE_74_io_sig_stat2trans)
  );
  PE PE_75 ( // @[pearray.scala 101:13]
    .clock(PE_75_clock),
    .reset(PE_75_reset),
    .io_data_2_in_bits(PE_75_io_data_2_in_bits),
    .io_data_2_out_bits(PE_75_io_data_2_out_bits),
    .io_data_1_in_valid(PE_75_io_data_1_in_valid),
    .io_data_1_in_bits(PE_75_io_data_1_in_bits),
    .io_data_1_out_valid(PE_75_io_data_1_out_valid),
    .io_data_1_out_bits(PE_75_io_data_1_out_bits),
    .io_data_0_in_valid(PE_75_io_data_0_in_valid),
    .io_data_0_in_bits(PE_75_io_data_0_in_bits),
    .io_data_0_out_valid(PE_75_io_data_0_out_valid),
    .io_data_0_out_bits(PE_75_io_data_0_out_bits),
    .io_sig_stat2trans(PE_75_io_sig_stat2trans)
  );
  PE PE_76 ( // @[pearray.scala 101:13]
    .clock(PE_76_clock),
    .reset(PE_76_reset),
    .io_data_2_in_bits(PE_76_io_data_2_in_bits),
    .io_data_2_out_bits(PE_76_io_data_2_out_bits),
    .io_data_1_in_valid(PE_76_io_data_1_in_valid),
    .io_data_1_in_bits(PE_76_io_data_1_in_bits),
    .io_data_1_out_valid(PE_76_io_data_1_out_valid),
    .io_data_1_out_bits(PE_76_io_data_1_out_bits),
    .io_data_0_in_valid(PE_76_io_data_0_in_valid),
    .io_data_0_in_bits(PE_76_io_data_0_in_bits),
    .io_data_0_out_valid(PE_76_io_data_0_out_valid),
    .io_data_0_out_bits(PE_76_io_data_0_out_bits),
    .io_sig_stat2trans(PE_76_io_sig_stat2trans)
  );
  PE PE_77 ( // @[pearray.scala 101:13]
    .clock(PE_77_clock),
    .reset(PE_77_reset),
    .io_data_2_in_bits(PE_77_io_data_2_in_bits),
    .io_data_2_out_bits(PE_77_io_data_2_out_bits),
    .io_data_1_in_valid(PE_77_io_data_1_in_valid),
    .io_data_1_in_bits(PE_77_io_data_1_in_bits),
    .io_data_1_out_valid(PE_77_io_data_1_out_valid),
    .io_data_1_out_bits(PE_77_io_data_1_out_bits),
    .io_data_0_in_valid(PE_77_io_data_0_in_valid),
    .io_data_0_in_bits(PE_77_io_data_0_in_bits),
    .io_data_0_out_valid(PE_77_io_data_0_out_valid),
    .io_data_0_out_bits(PE_77_io_data_0_out_bits),
    .io_sig_stat2trans(PE_77_io_sig_stat2trans)
  );
  PE PE_78 ( // @[pearray.scala 101:13]
    .clock(PE_78_clock),
    .reset(PE_78_reset),
    .io_data_2_in_bits(PE_78_io_data_2_in_bits),
    .io_data_2_out_bits(PE_78_io_data_2_out_bits),
    .io_data_1_in_valid(PE_78_io_data_1_in_valid),
    .io_data_1_in_bits(PE_78_io_data_1_in_bits),
    .io_data_1_out_valid(PE_78_io_data_1_out_valid),
    .io_data_1_out_bits(PE_78_io_data_1_out_bits),
    .io_data_0_in_valid(PE_78_io_data_0_in_valid),
    .io_data_0_in_bits(PE_78_io_data_0_in_bits),
    .io_data_0_out_valid(PE_78_io_data_0_out_valid),
    .io_data_0_out_bits(PE_78_io_data_0_out_bits),
    .io_sig_stat2trans(PE_78_io_sig_stat2trans)
  );
  PE PE_79 ( // @[pearray.scala 101:13]
    .clock(PE_79_clock),
    .reset(PE_79_reset),
    .io_data_2_in_bits(PE_79_io_data_2_in_bits),
    .io_data_2_out_bits(PE_79_io_data_2_out_bits),
    .io_data_1_in_valid(PE_79_io_data_1_in_valid),
    .io_data_1_in_bits(PE_79_io_data_1_in_bits),
    .io_data_1_out_valid(PE_79_io_data_1_out_valid),
    .io_data_1_out_bits(PE_79_io_data_1_out_bits),
    .io_data_0_in_valid(PE_79_io_data_0_in_valid),
    .io_data_0_in_bits(PE_79_io_data_0_in_bits),
    .io_data_0_out_valid(PE_79_io_data_0_out_valid),
    .io_data_0_out_bits(PE_79_io_data_0_out_bits),
    .io_sig_stat2trans(PE_79_io_sig_stat2trans)
  );
  PE PE_80 ( // @[pearray.scala 101:13]
    .clock(PE_80_clock),
    .reset(PE_80_reset),
    .io_data_2_in_bits(PE_80_io_data_2_in_bits),
    .io_data_2_out_bits(PE_80_io_data_2_out_bits),
    .io_data_1_in_valid(PE_80_io_data_1_in_valid),
    .io_data_1_in_bits(PE_80_io_data_1_in_bits),
    .io_data_1_out_valid(PE_80_io_data_1_out_valid),
    .io_data_1_out_bits(PE_80_io_data_1_out_bits),
    .io_data_0_in_valid(PE_80_io_data_0_in_valid),
    .io_data_0_in_bits(PE_80_io_data_0_in_bits),
    .io_data_0_out_valid(PE_80_io_data_0_out_valid),
    .io_data_0_out_bits(PE_80_io_data_0_out_bits),
    .io_sig_stat2trans(PE_80_io_sig_stat2trans)
  );
  PE PE_81 ( // @[pearray.scala 101:13]
    .clock(PE_81_clock),
    .reset(PE_81_reset),
    .io_data_2_in_bits(PE_81_io_data_2_in_bits),
    .io_data_2_out_bits(PE_81_io_data_2_out_bits),
    .io_data_1_in_valid(PE_81_io_data_1_in_valid),
    .io_data_1_in_bits(PE_81_io_data_1_in_bits),
    .io_data_1_out_valid(PE_81_io_data_1_out_valid),
    .io_data_1_out_bits(PE_81_io_data_1_out_bits),
    .io_data_0_in_valid(PE_81_io_data_0_in_valid),
    .io_data_0_in_bits(PE_81_io_data_0_in_bits),
    .io_data_0_out_valid(PE_81_io_data_0_out_valid),
    .io_data_0_out_bits(PE_81_io_data_0_out_bits),
    .io_sig_stat2trans(PE_81_io_sig_stat2trans)
  );
  PE PE_82 ( // @[pearray.scala 101:13]
    .clock(PE_82_clock),
    .reset(PE_82_reset),
    .io_data_2_in_bits(PE_82_io_data_2_in_bits),
    .io_data_2_out_bits(PE_82_io_data_2_out_bits),
    .io_data_1_in_valid(PE_82_io_data_1_in_valid),
    .io_data_1_in_bits(PE_82_io_data_1_in_bits),
    .io_data_1_out_valid(PE_82_io_data_1_out_valid),
    .io_data_1_out_bits(PE_82_io_data_1_out_bits),
    .io_data_0_in_valid(PE_82_io_data_0_in_valid),
    .io_data_0_in_bits(PE_82_io_data_0_in_bits),
    .io_data_0_out_valid(PE_82_io_data_0_out_valid),
    .io_data_0_out_bits(PE_82_io_data_0_out_bits),
    .io_sig_stat2trans(PE_82_io_sig_stat2trans)
  );
  PE PE_83 ( // @[pearray.scala 101:13]
    .clock(PE_83_clock),
    .reset(PE_83_reset),
    .io_data_2_in_bits(PE_83_io_data_2_in_bits),
    .io_data_2_out_bits(PE_83_io_data_2_out_bits),
    .io_data_1_in_valid(PE_83_io_data_1_in_valid),
    .io_data_1_in_bits(PE_83_io_data_1_in_bits),
    .io_data_1_out_valid(PE_83_io_data_1_out_valid),
    .io_data_1_out_bits(PE_83_io_data_1_out_bits),
    .io_data_0_in_valid(PE_83_io_data_0_in_valid),
    .io_data_0_in_bits(PE_83_io_data_0_in_bits),
    .io_data_0_out_valid(PE_83_io_data_0_out_valid),
    .io_data_0_out_bits(PE_83_io_data_0_out_bits),
    .io_sig_stat2trans(PE_83_io_sig_stat2trans)
  );
  PE PE_84 ( // @[pearray.scala 101:13]
    .clock(PE_84_clock),
    .reset(PE_84_reset),
    .io_data_2_in_bits(PE_84_io_data_2_in_bits),
    .io_data_2_out_bits(PE_84_io_data_2_out_bits),
    .io_data_1_in_valid(PE_84_io_data_1_in_valid),
    .io_data_1_in_bits(PE_84_io_data_1_in_bits),
    .io_data_1_out_valid(PE_84_io_data_1_out_valid),
    .io_data_1_out_bits(PE_84_io_data_1_out_bits),
    .io_data_0_in_valid(PE_84_io_data_0_in_valid),
    .io_data_0_in_bits(PE_84_io_data_0_in_bits),
    .io_data_0_out_valid(PE_84_io_data_0_out_valid),
    .io_data_0_out_bits(PE_84_io_data_0_out_bits),
    .io_sig_stat2trans(PE_84_io_sig_stat2trans)
  );
  PE PE_85 ( // @[pearray.scala 101:13]
    .clock(PE_85_clock),
    .reset(PE_85_reset),
    .io_data_2_in_bits(PE_85_io_data_2_in_bits),
    .io_data_2_out_bits(PE_85_io_data_2_out_bits),
    .io_data_1_in_valid(PE_85_io_data_1_in_valid),
    .io_data_1_in_bits(PE_85_io_data_1_in_bits),
    .io_data_1_out_valid(PE_85_io_data_1_out_valid),
    .io_data_1_out_bits(PE_85_io_data_1_out_bits),
    .io_data_0_in_valid(PE_85_io_data_0_in_valid),
    .io_data_0_in_bits(PE_85_io_data_0_in_bits),
    .io_data_0_out_valid(PE_85_io_data_0_out_valid),
    .io_data_0_out_bits(PE_85_io_data_0_out_bits),
    .io_sig_stat2trans(PE_85_io_sig_stat2trans)
  );
  PE PE_86 ( // @[pearray.scala 101:13]
    .clock(PE_86_clock),
    .reset(PE_86_reset),
    .io_data_2_in_bits(PE_86_io_data_2_in_bits),
    .io_data_2_out_bits(PE_86_io_data_2_out_bits),
    .io_data_1_in_valid(PE_86_io_data_1_in_valid),
    .io_data_1_in_bits(PE_86_io_data_1_in_bits),
    .io_data_1_out_valid(PE_86_io_data_1_out_valid),
    .io_data_1_out_bits(PE_86_io_data_1_out_bits),
    .io_data_0_in_valid(PE_86_io_data_0_in_valid),
    .io_data_0_in_bits(PE_86_io_data_0_in_bits),
    .io_data_0_out_valid(PE_86_io_data_0_out_valid),
    .io_data_0_out_bits(PE_86_io_data_0_out_bits),
    .io_sig_stat2trans(PE_86_io_sig_stat2trans)
  );
  PE PE_87 ( // @[pearray.scala 101:13]
    .clock(PE_87_clock),
    .reset(PE_87_reset),
    .io_data_2_in_bits(PE_87_io_data_2_in_bits),
    .io_data_2_out_bits(PE_87_io_data_2_out_bits),
    .io_data_1_in_valid(PE_87_io_data_1_in_valid),
    .io_data_1_in_bits(PE_87_io_data_1_in_bits),
    .io_data_1_out_valid(PE_87_io_data_1_out_valid),
    .io_data_1_out_bits(PE_87_io_data_1_out_bits),
    .io_data_0_in_valid(PE_87_io_data_0_in_valid),
    .io_data_0_in_bits(PE_87_io_data_0_in_bits),
    .io_data_0_out_valid(PE_87_io_data_0_out_valid),
    .io_data_0_out_bits(PE_87_io_data_0_out_bits),
    .io_sig_stat2trans(PE_87_io_sig_stat2trans)
  );
  PE PE_88 ( // @[pearray.scala 101:13]
    .clock(PE_88_clock),
    .reset(PE_88_reset),
    .io_data_2_in_bits(PE_88_io_data_2_in_bits),
    .io_data_2_out_bits(PE_88_io_data_2_out_bits),
    .io_data_1_in_valid(PE_88_io_data_1_in_valid),
    .io_data_1_in_bits(PE_88_io_data_1_in_bits),
    .io_data_1_out_valid(PE_88_io_data_1_out_valid),
    .io_data_1_out_bits(PE_88_io_data_1_out_bits),
    .io_data_0_in_valid(PE_88_io_data_0_in_valid),
    .io_data_0_in_bits(PE_88_io_data_0_in_bits),
    .io_data_0_out_valid(PE_88_io_data_0_out_valid),
    .io_data_0_out_bits(PE_88_io_data_0_out_bits),
    .io_sig_stat2trans(PE_88_io_sig_stat2trans)
  );
  PE PE_89 ( // @[pearray.scala 101:13]
    .clock(PE_89_clock),
    .reset(PE_89_reset),
    .io_data_2_in_bits(PE_89_io_data_2_in_bits),
    .io_data_2_out_bits(PE_89_io_data_2_out_bits),
    .io_data_1_in_valid(PE_89_io_data_1_in_valid),
    .io_data_1_in_bits(PE_89_io_data_1_in_bits),
    .io_data_1_out_valid(PE_89_io_data_1_out_valid),
    .io_data_1_out_bits(PE_89_io_data_1_out_bits),
    .io_data_0_in_valid(PE_89_io_data_0_in_valid),
    .io_data_0_in_bits(PE_89_io_data_0_in_bits),
    .io_data_0_out_valid(PE_89_io_data_0_out_valid),
    .io_data_0_out_bits(PE_89_io_data_0_out_bits),
    .io_sig_stat2trans(PE_89_io_sig_stat2trans)
  );
  PE PE_90 ( // @[pearray.scala 101:13]
    .clock(PE_90_clock),
    .reset(PE_90_reset),
    .io_data_2_in_bits(PE_90_io_data_2_in_bits),
    .io_data_2_out_bits(PE_90_io_data_2_out_bits),
    .io_data_1_in_valid(PE_90_io_data_1_in_valid),
    .io_data_1_in_bits(PE_90_io_data_1_in_bits),
    .io_data_1_out_valid(PE_90_io_data_1_out_valid),
    .io_data_1_out_bits(PE_90_io_data_1_out_bits),
    .io_data_0_in_valid(PE_90_io_data_0_in_valid),
    .io_data_0_in_bits(PE_90_io_data_0_in_bits),
    .io_data_0_out_valid(PE_90_io_data_0_out_valid),
    .io_data_0_out_bits(PE_90_io_data_0_out_bits),
    .io_sig_stat2trans(PE_90_io_sig_stat2trans)
  );
  PE PE_91 ( // @[pearray.scala 101:13]
    .clock(PE_91_clock),
    .reset(PE_91_reset),
    .io_data_2_in_bits(PE_91_io_data_2_in_bits),
    .io_data_2_out_bits(PE_91_io_data_2_out_bits),
    .io_data_1_in_valid(PE_91_io_data_1_in_valid),
    .io_data_1_in_bits(PE_91_io_data_1_in_bits),
    .io_data_1_out_valid(PE_91_io_data_1_out_valid),
    .io_data_1_out_bits(PE_91_io_data_1_out_bits),
    .io_data_0_in_valid(PE_91_io_data_0_in_valid),
    .io_data_0_in_bits(PE_91_io_data_0_in_bits),
    .io_data_0_out_valid(PE_91_io_data_0_out_valid),
    .io_data_0_out_bits(PE_91_io_data_0_out_bits),
    .io_sig_stat2trans(PE_91_io_sig_stat2trans)
  );
  PE PE_92 ( // @[pearray.scala 101:13]
    .clock(PE_92_clock),
    .reset(PE_92_reset),
    .io_data_2_in_bits(PE_92_io_data_2_in_bits),
    .io_data_2_out_bits(PE_92_io_data_2_out_bits),
    .io_data_1_in_valid(PE_92_io_data_1_in_valid),
    .io_data_1_in_bits(PE_92_io_data_1_in_bits),
    .io_data_1_out_valid(PE_92_io_data_1_out_valid),
    .io_data_1_out_bits(PE_92_io_data_1_out_bits),
    .io_data_0_in_valid(PE_92_io_data_0_in_valid),
    .io_data_0_in_bits(PE_92_io_data_0_in_bits),
    .io_data_0_out_valid(PE_92_io_data_0_out_valid),
    .io_data_0_out_bits(PE_92_io_data_0_out_bits),
    .io_sig_stat2trans(PE_92_io_sig_stat2trans)
  );
  PE PE_93 ( // @[pearray.scala 101:13]
    .clock(PE_93_clock),
    .reset(PE_93_reset),
    .io_data_2_in_bits(PE_93_io_data_2_in_bits),
    .io_data_2_out_bits(PE_93_io_data_2_out_bits),
    .io_data_1_in_valid(PE_93_io_data_1_in_valid),
    .io_data_1_in_bits(PE_93_io_data_1_in_bits),
    .io_data_1_out_valid(PE_93_io_data_1_out_valid),
    .io_data_1_out_bits(PE_93_io_data_1_out_bits),
    .io_data_0_in_valid(PE_93_io_data_0_in_valid),
    .io_data_0_in_bits(PE_93_io_data_0_in_bits),
    .io_data_0_out_valid(PE_93_io_data_0_out_valid),
    .io_data_0_out_bits(PE_93_io_data_0_out_bits),
    .io_sig_stat2trans(PE_93_io_sig_stat2trans)
  );
  PE PE_94 ( // @[pearray.scala 101:13]
    .clock(PE_94_clock),
    .reset(PE_94_reset),
    .io_data_2_in_bits(PE_94_io_data_2_in_bits),
    .io_data_2_out_bits(PE_94_io_data_2_out_bits),
    .io_data_1_in_valid(PE_94_io_data_1_in_valid),
    .io_data_1_in_bits(PE_94_io_data_1_in_bits),
    .io_data_1_out_valid(PE_94_io_data_1_out_valid),
    .io_data_1_out_bits(PE_94_io_data_1_out_bits),
    .io_data_0_in_valid(PE_94_io_data_0_in_valid),
    .io_data_0_in_bits(PE_94_io_data_0_in_bits),
    .io_data_0_out_valid(PE_94_io_data_0_out_valid),
    .io_data_0_out_bits(PE_94_io_data_0_out_bits),
    .io_sig_stat2trans(PE_94_io_sig_stat2trans)
  );
  PE PE_95 ( // @[pearray.scala 101:13]
    .clock(PE_95_clock),
    .reset(PE_95_reset),
    .io_data_2_in_bits(PE_95_io_data_2_in_bits),
    .io_data_2_out_bits(PE_95_io_data_2_out_bits),
    .io_data_1_in_valid(PE_95_io_data_1_in_valid),
    .io_data_1_in_bits(PE_95_io_data_1_in_bits),
    .io_data_1_out_valid(PE_95_io_data_1_out_valid),
    .io_data_1_out_bits(PE_95_io_data_1_out_bits),
    .io_data_0_in_valid(PE_95_io_data_0_in_valid),
    .io_data_0_in_bits(PE_95_io_data_0_in_bits),
    .io_data_0_out_valid(PE_95_io_data_0_out_valid),
    .io_data_0_out_bits(PE_95_io_data_0_out_bits),
    .io_sig_stat2trans(PE_95_io_sig_stat2trans)
  );
  PE PE_96 ( // @[pearray.scala 101:13]
    .clock(PE_96_clock),
    .reset(PE_96_reset),
    .io_data_2_in_bits(PE_96_io_data_2_in_bits),
    .io_data_2_out_bits(PE_96_io_data_2_out_bits),
    .io_data_1_in_valid(PE_96_io_data_1_in_valid),
    .io_data_1_in_bits(PE_96_io_data_1_in_bits),
    .io_data_1_out_valid(PE_96_io_data_1_out_valid),
    .io_data_1_out_bits(PE_96_io_data_1_out_bits),
    .io_data_0_in_valid(PE_96_io_data_0_in_valid),
    .io_data_0_in_bits(PE_96_io_data_0_in_bits),
    .io_data_0_out_valid(PE_96_io_data_0_out_valid),
    .io_data_0_out_bits(PE_96_io_data_0_out_bits),
    .io_sig_stat2trans(PE_96_io_sig_stat2trans)
  );
  PE PE_97 ( // @[pearray.scala 101:13]
    .clock(PE_97_clock),
    .reset(PE_97_reset),
    .io_data_2_in_bits(PE_97_io_data_2_in_bits),
    .io_data_2_out_bits(PE_97_io_data_2_out_bits),
    .io_data_1_in_valid(PE_97_io_data_1_in_valid),
    .io_data_1_in_bits(PE_97_io_data_1_in_bits),
    .io_data_1_out_valid(PE_97_io_data_1_out_valid),
    .io_data_1_out_bits(PE_97_io_data_1_out_bits),
    .io_data_0_in_valid(PE_97_io_data_0_in_valid),
    .io_data_0_in_bits(PE_97_io_data_0_in_bits),
    .io_data_0_out_valid(PE_97_io_data_0_out_valid),
    .io_data_0_out_bits(PE_97_io_data_0_out_bits),
    .io_sig_stat2trans(PE_97_io_sig_stat2trans)
  );
  PE PE_98 ( // @[pearray.scala 101:13]
    .clock(PE_98_clock),
    .reset(PE_98_reset),
    .io_data_2_in_bits(PE_98_io_data_2_in_bits),
    .io_data_2_out_bits(PE_98_io_data_2_out_bits),
    .io_data_1_in_valid(PE_98_io_data_1_in_valid),
    .io_data_1_in_bits(PE_98_io_data_1_in_bits),
    .io_data_1_out_valid(PE_98_io_data_1_out_valid),
    .io_data_1_out_bits(PE_98_io_data_1_out_bits),
    .io_data_0_in_valid(PE_98_io_data_0_in_valid),
    .io_data_0_in_bits(PE_98_io_data_0_in_bits),
    .io_data_0_out_valid(PE_98_io_data_0_out_valid),
    .io_data_0_out_bits(PE_98_io_data_0_out_bits),
    .io_sig_stat2trans(PE_98_io_sig_stat2trans)
  );
  PE PE_99 ( // @[pearray.scala 101:13]
    .clock(PE_99_clock),
    .reset(PE_99_reset),
    .io_data_2_in_bits(PE_99_io_data_2_in_bits),
    .io_data_2_out_bits(PE_99_io_data_2_out_bits),
    .io_data_1_in_valid(PE_99_io_data_1_in_valid),
    .io_data_1_in_bits(PE_99_io_data_1_in_bits),
    .io_data_1_out_valid(PE_99_io_data_1_out_valid),
    .io_data_1_out_bits(PE_99_io_data_1_out_bits),
    .io_data_0_in_valid(PE_99_io_data_0_in_valid),
    .io_data_0_in_bits(PE_99_io_data_0_in_bits),
    .io_data_0_out_valid(PE_99_io_data_0_out_valid),
    .io_data_0_out_bits(PE_99_io_data_0_out_bits),
    .io_sig_stat2trans(PE_99_io_sig_stat2trans)
  );
  PE PE_100 ( // @[pearray.scala 101:13]
    .clock(PE_100_clock),
    .reset(PE_100_reset),
    .io_data_2_in_bits(PE_100_io_data_2_in_bits),
    .io_data_2_out_bits(PE_100_io_data_2_out_bits),
    .io_data_1_in_valid(PE_100_io_data_1_in_valid),
    .io_data_1_in_bits(PE_100_io_data_1_in_bits),
    .io_data_1_out_valid(PE_100_io_data_1_out_valid),
    .io_data_1_out_bits(PE_100_io_data_1_out_bits),
    .io_data_0_in_valid(PE_100_io_data_0_in_valid),
    .io_data_0_in_bits(PE_100_io_data_0_in_bits),
    .io_data_0_out_valid(PE_100_io_data_0_out_valid),
    .io_data_0_out_bits(PE_100_io_data_0_out_bits),
    .io_sig_stat2trans(PE_100_io_sig_stat2trans)
  );
  PE PE_101 ( // @[pearray.scala 101:13]
    .clock(PE_101_clock),
    .reset(PE_101_reset),
    .io_data_2_in_bits(PE_101_io_data_2_in_bits),
    .io_data_2_out_bits(PE_101_io_data_2_out_bits),
    .io_data_1_in_valid(PE_101_io_data_1_in_valid),
    .io_data_1_in_bits(PE_101_io_data_1_in_bits),
    .io_data_1_out_valid(PE_101_io_data_1_out_valid),
    .io_data_1_out_bits(PE_101_io_data_1_out_bits),
    .io_data_0_in_valid(PE_101_io_data_0_in_valid),
    .io_data_0_in_bits(PE_101_io_data_0_in_bits),
    .io_data_0_out_valid(PE_101_io_data_0_out_valid),
    .io_data_0_out_bits(PE_101_io_data_0_out_bits),
    .io_sig_stat2trans(PE_101_io_sig_stat2trans)
  );
  PE PE_102 ( // @[pearray.scala 101:13]
    .clock(PE_102_clock),
    .reset(PE_102_reset),
    .io_data_2_in_bits(PE_102_io_data_2_in_bits),
    .io_data_2_out_bits(PE_102_io_data_2_out_bits),
    .io_data_1_in_valid(PE_102_io_data_1_in_valid),
    .io_data_1_in_bits(PE_102_io_data_1_in_bits),
    .io_data_1_out_valid(PE_102_io_data_1_out_valid),
    .io_data_1_out_bits(PE_102_io_data_1_out_bits),
    .io_data_0_in_valid(PE_102_io_data_0_in_valid),
    .io_data_0_in_bits(PE_102_io_data_0_in_bits),
    .io_data_0_out_valid(PE_102_io_data_0_out_valid),
    .io_data_0_out_bits(PE_102_io_data_0_out_bits),
    .io_sig_stat2trans(PE_102_io_sig_stat2trans)
  );
  PE PE_103 ( // @[pearray.scala 101:13]
    .clock(PE_103_clock),
    .reset(PE_103_reset),
    .io_data_2_in_bits(PE_103_io_data_2_in_bits),
    .io_data_2_out_bits(PE_103_io_data_2_out_bits),
    .io_data_1_in_valid(PE_103_io_data_1_in_valid),
    .io_data_1_in_bits(PE_103_io_data_1_in_bits),
    .io_data_1_out_valid(PE_103_io_data_1_out_valid),
    .io_data_1_out_bits(PE_103_io_data_1_out_bits),
    .io_data_0_in_valid(PE_103_io_data_0_in_valid),
    .io_data_0_in_bits(PE_103_io_data_0_in_bits),
    .io_data_0_out_valid(PE_103_io_data_0_out_valid),
    .io_data_0_out_bits(PE_103_io_data_0_out_bits),
    .io_sig_stat2trans(PE_103_io_sig_stat2trans)
  );
  PE PE_104 ( // @[pearray.scala 101:13]
    .clock(PE_104_clock),
    .reset(PE_104_reset),
    .io_data_2_in_bits(PE_104_io_data_2_in_bits),
    .io_data_2_out_bits(PE_104_io_data_2_out_bits),
    .io_data_1_in_valid(PE_104_io_data_1_in_valid),
    .io_data_1_in_bits(PE_104_io_data_1_in_bits),
    .io_data_1_out_valid(PE_104_io_data_1_out_valid),
    .io_data_1_out_bits(PE_104_io_data_1_out_bits),
    .io_data_0_in_valid(PE_104_io_data_0_in_valid),
    .io_data_0_in_bits(PE_104_io_data_0_in_bits),
    .io_data_0_out_valid(PE_104_io_data_0_out_valid),
    .io_data_0_out_bits(PE_104_io_data_0_out_bits),
    .io_sig_stat2trans(PE_104_io_sig_stat2trans)
  );
  PE PE_105 ( // @[pearray.scala 101:13]
    .clock(PE_105_clock),
    .reset(PE_105_reset),
    .io_data_2_in_bits(PE_105_io_data_2_in_bits),
    .io_data_2_out_bits(PE_105_io_data_2_out_bits),
    .io_data_1_in_valid(PE_105_io_data_1_in_valid),
    .io_data_1_in_bits(PE_105_io_data_1_in_bits),
    .io_data_1_out_valid(PE_105_io_data_1_out_valid),
    .io_data_1_out_bits(PE_105_io_data_1_out_bits),
    .io_data_0_in_valid(PE_105_io_data_0_in_valid),
    .io_data_0_in_bits(PE_105_io_data_0_in_bits),
    .io_data_0_out_valid(PE_105_io_data_0_out_valid),
    .io_data_0_out_bits(PE_105_io_data_0_out_bits),
    .io_sig_stat2trans(PE_105_io_sig_stat2trans)
  );
  PE PE_106 ( // @[pearray.scala 101:13]
    .clock(PE_106_clock),
    .reset(PE_106_reset),
    .io_data_2_in_bits(PE_106_io_data_2_in_bits),
    .io_data_2_out_bits(PE_106_io_data_2_out_bits),
    .io_data_1_in_valid(PE_106_io_data_1_in_valid),
    .io_data_1_in_bits(PE_106_io_data_1_in_bits),
    .io_data_1_out_valid(PE_106_io_data_1_out_valid),
    .io_data_1_out_bits(PE_106_io_data_1_out_bits),
    .io_data_0_in_valid(PE_106_io_data_0_in_valid),
    .io_data_0_in_bits(PE_106_io_data_0_in_bits),
    .io_data_0_out_valid(PE_106_io_data_0_out_valid),
    .io_data_0_out_bits(PE_106_io_data_0_out_bits),
    .io_sig_stat2trans(PE_106_io_sig_stat2trans)
  );
  PE PE_107 ( // @[pearray.scala 101:13]
    .clock(PE_107_clock),
    .reset(PE_107_reset),
    .io_data_2_in_bits(PE_107_io_data_2_in_bits),
    .io_data_2_out_bits(PE_107_io_data_2_out_bits),
    .io_data_1_in_valid(PE_107_io_data_1_in_valid),
    .io_data_1_in_bits(PE_107_io_data_1_in_bits),
    .io_data_1_out_valid(PE_107_io_data_1_out_valid),
    .io_data_1_out_bits(PE_107_io_data_1_out_bits),
    .io_data_0_in_valid(PE_107_io_data_0_in_valid),
    .io_data_0_in_bits(PE_107_io_data_0_in_bits),
    .io_data_0_out_valid(PE_107_io_data_0_out_valid),
    .io_data_0_out_bits(PE_107_io_data_0_out_bits),
    .io_sig_stat2trans(PE_107_io_sig_stat2trans)
  );
  PE PE_108 ( // @[pearray.scala 101:13]
    .clock(PE_108_clock),
    .reset(PE_108_reset),
    .io_data_2_in_bits(PE_108_io_data_2_in_bits),
    .io_data_2_out_bits(PE_108_io_data_2_out_bits),
    .io_data_1_in_valid(PE_108_io_data_1_in_valid),
    .io_data_1_in_bits(PE_108_io_data_1_in_bits),
    .io_data_1_out_valid(PE_108_io_data_1_out_valid),
    .io_data_1_out_bits(PE_108_io_data_1_out_bits),
    .io_data_0_in_valid(PE_108_io_data_0_in_valid),
    .io_data_0_in_bits(PE_108_io_data_0_in_bits),
    .io_data_0_out_valid(PE_108_io_data_0_out_valid),
    .io_data_0_out_bits(PE_108_io_data_0_out_bits),
    .io_sig_stat2trans(PE_108_io_sig_stat2trans)
  );
  PE PE_109 ( // @[pearray.scala 101:13]
    .clock(PE_109_clock),
    .reset(PE_109_reset),
    .io_data_2_in_bits(PE_109_io_data_2_in_bits),
    .io_data_2_out_bits(PE_109_io_data_2_out_bits),
    .io_data_1_in_valid(PE_109_io_data_1_in_valid),
    .io_data_1_in_bits(PE_109_io_data_1_in_bits),
    .io_data_1_out_valid(PE_109_io_data_1_out_valid),
    .io_data_1_out_bits(PE_109_io_data_1_out_bits),
    .io_data_0_in_valid(PE_109_io_data_0_in_valid),
    .io_data_0_in_bits(PE_109_io_data_0_in_bits),
    .io_data_0_out_valid(PE_109_io_data_0_out_valid),
    .io_data_0_out_bits(PE_109_io_data_0_out_bits),
    .io_sig_stat2trans(PE_109_io_sig_stat2trans)
  );
  PE PE_110 ( // @[pearray.scala 101:13]
    .clock(PE_110_clock),
    .reset(PE_110_reset),
    .io_data_2_in_bits(PE_110_io_data_2_in_bits),
    .io_data_2_out_bits(PE_110_io_data_2_out_bits),
    .io_data_1_in_valid(PE_110_io_data_1_in_valid),
    .io_data_1_in_bits(PE_110_io_data_1_in_bits),
    .io_data_1_out_valid(PE_110_io_data_1_out_valid),
    .io_data_1_out_bits(PE_110_io_data_1_out_bits),
    .io_data_0_in_valid(PE_110_io_data_0_in_valid),
    .io_data_0_in_bits(PE_110_io_data_0_in_bits),
    .io_data_0_out_valid(PE_110_io_data_0_out_valid),
    .io_data_0_out_bits(PE_110_io_data_0_out_bits),
    .io_sig_stat2trans(PE_110_io_sig_stat2trans)
  );
  PE PE_111 ( // @[pearray.scala 101:13]
    .clock(PE_111_clock),
    .reset(PE_111_reset),
    .io_data_2_in_bits(PE_111_io_data_2_in_bits),
    .io_data_2_out_bits(PE_111_io_data_2_out_bits),
    .io_data_1_in_valid(PE_111_io_data_1_in_valid),
    .io_data_1_in_bits(PE_111_io_data_1_in_bits),
    .io_data_1_out_valid(PE_111_io_data_1_out_valid),
    .io_data_1_out_bits(PE_111_io_data_1_out_bits),
    .io_data_0_in_valid(PE_111_io_data_0_in_valid),
    .io_data_0_in_bits(PE_111_io_data_0_in_bits),
    .io_data_0_out_valid(PE_111_io_data_0_out_valid),
    .io_data_0_out_bits(PE_111_io_data_0_out_bits),
    .io_sig_stat2trans(PE_111_io_sig_stat2trans)
  );
  PE PE_112 ( // @[pearray.scala 101:13]
    .clock(PE_112_clock),
    .reset(PE_112_reset),
    .io_data_2_in_bits(PE_112_io_data_2_in_bits),
    .io_data_2_out_bits(PE_112_io_data_2_out_bits),
    .io_data_1_in_valid(PE_112_io_data_1_in_valid),
    .io_data_1_in_bits(PE_112_io_data_1_in_bits),
    .io_data_1_out_valid(PE_112_io_data_1_out_valid),
    .io_data_1_out_bits(PE_112_io_data_1_out_bits),
    .io_data_0_in_valid(PE_112_io_data_0_in_valid),
    .io_data_0_in_bits(PE_112_io_data_0_in_bits),
    .io_data_0_out_valid(PE_112_io_data_0_out_valid),
    .io_data_0_out_bits(PE_112_io_data_0_out_bits),
    .io_sig_stat2trans(PE_112_io_sig_stat2trans)
  );
  PE PE_113 ( // @[pearray.scala 101:13]
    .clock(PE_113_clock),
    .reset(PE_113_reset),
    .io_data_2_in_bits(PE_113_io_data_2_in_bits),
    .io_data_2_out_bits(PE_113_io_data_2_out_bits),
    .io_data_1_in_valid(PE_113_io_data_1_in_valid),
    .io_data_1_in_bits(PE_113_io_data_1_in_bits),
    .io_data_1_out_valid(PE_113_io_data_1_out_valid),
    .io_data_1_out_bits(PE_113_io_data_1_out_bits),
    .io_data_0_in_valid(PE_113_io_data_0_in_valid),
    .io_data_0_in_bits(PE_113_io_data_0_in_bits),
    .io_data_0_out_valid(PE_113_io_data_0_out_valid),
    .io_data_0_out_bits(PE_113_io_data_0_out_bits),
    .io_sig_stat2trans(PE_113_io_sig_stat2trans)
  );
  PE PE_114 ( // @[pearray.scala 101:13]
    .clock(PE_114_clock),
    .reset(PE_114_reset),
    .io_data_2_in_bits(PE_114_io_data_2_in_bits),
    .io_data_2_out_bits(PE_114_io_data_2_out_bits),
    .io_data_1_in_valid(PE_114_io_data_1_in_valid),
    .io_data_1_in_bits(PE_114_io_data_1_in_bits),
    .io_data_1_out_valid(PE_114_io_data_1_out_valid),
    .io_data_1_out_bits(PE_114_io_data_1_out_bits),
    .io_data_0_in_valid(PE_114_io_data_0_in_valid),
    .io_data_0_in_bits(PE_114_io_data_0_in_bits),
    .io_data_0_out_valid(PE_114_io_data_0_out_valid),
    .io_data_0_out_bits(PE_114_io_data_0_out_bits),
    .io_sig_stat2trans(PE_114_io_sig_stat2trans)
  );
  PE PE_115 ( // @[pearray.scala 101:13]
    .clock(PE_115_clock),
    .reset(PE_115_reset),
    .io_data_2_in_bits(PE_115_io_data_2_in_bits),
    .io_data_2_out_bits(PE_115_io_data_2_out_bits),
    .io_data_1_in_valid(PE_115_io_data_1_in_valid),
    .io_data_1_in_bits(PE_115_io_data_1_in_bits),
    .io_data_1_out_valid(PE_115_io_data_1_out_valid),
    .io_data_1_out_bits(PE_115_io_data_1_out_bits),
    .io_data_0_in_valid(PE_115_io_data_0_in_valid),
    .io_data_0_in_bits(PE_115_io_data_0_in_bits),
    .io_data_0_out_valid(PE_115_io_data_0_out_valid),
    .io_data_0_out_bits(PE_115_io_data_0_out_bits),
    .io_sig_stat2trans(PE_115_io_sig_stat2trans)
  );
  PE PE_116 ( // @[pearray.scala 101:13]
    .clock(PE_116_clock),
    .reset(PE_116_reset),
    .io_data_2_in_bits(PE_116_io_data_2_in_bits),
    .io_data_2_out_bits(PE_116_io_data_2_out_bits),
    .io_data_1_in_valid(PE_116_io_data_1_in_valid),
    .io_data_1_in_bits(PE_116_io_data_1_in_bits),
    .io_data_1_out_valid(PE_116_io_data_1_out_valid),
    .io_data_1_out_bits(PE_116_io_data_1_out_bits),
    .io_data_0_in_valid(PE_116_io_data_0_in_valid),
    .io_data_0_in_bits(PE_116_io_data_0_in_bits),
    .io_data_0_out_valid(PE_116_io_data_0_out_valid),
    .io_data_0_out_bits(PE_116_io_data_0_out_bits),
    .io_sig_stat2trans(PE_116_io_sig_stat2trans)
  );
  PE PE_117 ( // @[pearray.scala 101:13]
    .clock(PE_117_clock),
    .reset(PE_117_reset),
    .io_data_2_in_bits(PE_117_io_data_2_in_bits),
    .io_data_2_out_bits(PE_117_io_data_2_out_bits),
    .io_data_1_in_valid(PE_117_io_data_1_in_valid),
    .io_data_1_in_bits(PE_117_io_data_1_in_bits),
    .io_data_1_out_valid(PE_117_io_data_1_out_valid),
    .io_data_1_out_bits(PE_117_io_data_1_out_bits),
    .io_data_0_in_valid(PE_117_io_data_0_in_valid),
    .io_data_0_in_bits(PE_117_io_data_0_in_bits),
    .io_data_0_out_valid(PE_117_io_data_0_out_valid),
    .io_data_0_out_bits(PE_117_io_data_0_out_bits),
    .io_sig_stat2trans(PE_117_io_sig_stat2trans)
  );
  PE PE_118 ( // @[pearray.scala 101:13]
    .clock(PE_118_clock),
    .reset(PE_118_reset),
    .io_data_2_in_bits(PE_118_io_data_2_in_bits),
    .io_data_2_out_bits(PE_118_io_data_2_out_bits),
    .io_data_1_in_valid(PE_118_io_data_1_in_valid),
    .io_data_1_in_bits(PE_118_io_data_1_in_bits),
    .io_data_1_out_valid(PE_118_io_data_1_out_valid),
    .io_data_1_out_bits(PE_118_io_data_1_out_bits),
    .io_data_0_in_valid(PE_118_io_data_0_in_valid),
    .io_data_0_in_bits(PE_118_io_data_0_in_bits),
    .io_data_0_out_valid(PE_118_io_data_0_out_valid),
    .io_data_0_out_bits(PE_118_io_data_0_out_bits),
    .io_sig_stat2trans(PE_118_io_sig_stat2trans)
  );
  PE PE_119 ( // @[pearray.scala 101:13]
    .clock(PE_119_clock),
    .reset(PE_119_reset),
    .io_data_2_in_bits(PE_119_io_data_2_in_bits),
    .io_data_2_out_bits(PE_119_io_data_2_out_bits),
    .io_data_1_in_valid(PE_119_io_data_1_in_valid),
    .io_data_1_in_bits(PE_119_io_data_1_in_bits),
    .io_data_1_out_valid(PE_119_io_data_1_out_valid),
    .io_data_1_out_bits(PE_119_io_data_1_out_bits),
    .io_data_0_in_valid(PE_119_io_data_0_in_valid),
    .io_data_0_in_bits(PE_119_io_data_0_in_bits),
    .io_data_0_out_valid(PE_119_io_data_0_out_valid),
    .io_data_0_out_bits(PE_119_io_data_0_out_bits),
    .io_sig_stat2trans(PE_119_io_sig_stat2trans)
  );
  PE PE_120 ( // @[pearray.scala 101:13]
    .clock(PE_120_clock),
    .reset(PE_120_reset),
    .io_data_2_in_bits(PE_120_io_data_2_in_bits),
    .io_data_2_out_bits(PE_120_io_data_2_out_bits),
    .io_data_1_in_valid(PE_120_io_data_1_in_valid),
    .io_data_1_in_bits(PE_120_io_data_1_in_bits),
    .io_data_1_out_valid(PE_120_io_data_1_out_valid),
    .io_data_1_out_bits(PE_120_io_data_1_out_bits),
    .io_data_0_in_valid(PE_120_io_data_0_in_valid),
    .io_data_0_in_bits(PE_120_io_data_0_in_bits),
    .io_data_0_out_valid(PE_120_io_data_0_out_valid),
    .io_data_0_out_bits(PE_120_io_data_0_out_bits),
    .io_sig_stat2trans(PE_120_io_sig_stat2trans)
  );
  PE PE_121 ( // @[pearray.scala 101:13]
    .clock(PE_121_clock),
    .reset(PE_121_reset),
    .io_data_2_in_bits(PE_121_io_data_2_in_bits),
    .io_data_2_out_bits(PE_121_io_data_2_out_bits),
    .io_data_1_in_valid(PE_121_io_data_1_in_valid),
    .io_data_1_in_bits(PE_121_io_data_1_in_bits),
    .io_data_1_out_valid(PE_121_io_data_1_out_valid),
    .io_data_1_out_bits(PE_121_io_data_1_out_bits),
    .io_data_0_in_valid(PE_121_io_data_0_in_valid),
    .io_data_0_in_bits(PE_121_io_data_0_in_bits),
    .io_data_0_out_valid(PE_121_io_data_0_out_valid),
    .io_data_0_out_bits(PE_121_io_data_0_out_bits),
    .io_sig_stat2trans(PE_121_io_sig_stat2trans)
  );
  PE PE_122 ( // @[pearray.scala 101:13]
    .clock(PE_122_clock),
    .reset(PE_122_reset),
    .io_data_2_in_bits(PE_122_io_data_2_in_bits),
    .io_data_2_out_bits(PE_122_io_data_2_out_bits),
    .io_data_1_in_valid(PE_122_io_data_1_in_valid),
    .io_data_1_in_bits(PE_122_io_data_1_in_bits),
    .io_data_1_out_valid(PE_122_io_data_1_out_valid),
    .io_data_1_out_bits(PE_122_io_data_1_out_bits),
    .io_data_0_in_valid(PE_122_io_data_0_in_valid),
    .io_data_0_in_bits(PE_122_io_data_0_in_bits),
    .io_data_0_out_valid(PE_122_io_data_0_out_valid),
    .io_data_0_out_bits(PE_122_io_data_0_out_bits),
    .io_sig_stat2trans(PE_122_io_sig_stat2trans)
  );
  PE PE_123 ( // @[pearray.scala 101:13]
    .clock(PE_123_clock),
    .reset(PE_123_reset),
    .io_data_2_in_bits(PE_123_io_data_2_in_bits),
    .io_data_2_out_bits(PE_123_io_data_2_out_bits),
    .io_data_1_in_valid(PE_123_io_data_1_in_valid),
    .io_data_1_in_bits(PE_123_io_data_1_in_bits),
    .io_data_1_out_valid(PE_123_io_data_1_out_valid),
    .io_data_1_out_bits(PE_123_io_data_1_out_bits),
    .io_data_0_in_valid(PE_123_io_data_0_in_valid),
    .io_data_0_in_bits(PE_123_io_data_0_in_bits),
    .io_data_0_out_valid(PE_123_io_data_0_out_valid),
    .io_data_0_out_bits(PE_123_io_data_0_out_bits),
    .io_sig_stat2trans(PE_123_io_sig_stat2trans)
  );
  PE PE_124 ( // @[pearray.scala 101:13]
    .clock(PE_124_clock),
    .reset(PE_124_reset),
    .io_data_2_in_bits(PE_124_io_data_2_in_bits),
    .io_data_2_out_bits(PE_124_io_data_2_out_bits),
    .io_data_1_in_valid(PE_124_io_data_1_in_valid),
    .io_data_1_in_bits(PE_124_io_data_1_in_bits),
    .io_data_1_out_valid(PE_124_io_data_1_out_valid),
    .io_data_1_out_bits(PE_124_io_data_1_out_bits),
    .io_data_0_in_valid(PE_124_io_data_0_in_valid),
    .io_data_0_in_bits(PE_124_io_data_0_in_bits),
    .io_data_0_out_valid(PE_124_io_data_0_out_valid),
    .io_data_0_out_bits(PE_124_io_data_0_out_bits),
    .io_sig_stat2trans(PE_124_io_sig_stat2trans)
  );
  PE PE_125 ( // @[pearray.scala 101:13]
    .clock(PE_125_clock),
    .reset(PE_125_reset),
    .io_data_2_in_bits(PE_125_io_data_2_in_bits),
    .io_data_2_out_bits(PE_125_io_data_2_out_bits),
    .io_data_1_in_valid(PE_125_io_data_1_in_valid),
    .io_data_1_in_bits(PE_125_io_data_1_in_bits),
    .io_data_1_out_valid(PE_125_io_data_1_out_valid),
    .io_data_1_out_bits(PE_125_io_data_1_out_bits),
    .io_data_0_in_valid(PE_125_io_data_0_in_valid),
    .io_data_0_in_bits(PE_125_io_data_0_in_bits),
    .io_data_0_out_valid(PE_125_io_data_0_out_valid),
    .io_data_0_out_bits(PE_125_io_data_0_out_bits),
    .io_sig_stat2trans(PE_125_io_sig_stat2trans)
  );
  PE PE_126 ( // @[pearray.scala 101:13]
    .clock(PE_126_clock),
    .reset(PE_126_reset),
    .io_data_2_in_bits(PE_126_io_data_2_in_bits),
    .io_data_2_out_bits(PE_126_io_data_2_out_bits),
    .io_data_1_in_valid(PE_126_io_data_1_in_valid),
    .io_data_1_in_bits(PE_126_io_data_1_in_bits),
    .io_data_1_out_valid(PE_126_io_data_1_out_valid),
    .io_data_1_out_bits(PE_126_io_data_1_out_bits),
    .io_data_0_in_valid(PE_126_io_data_0_in_valid),
    .io_data_0_in_bits(PE_126_io_data_0_in_bits),
    .io_data_0_out_valid(PE_126_io_data_0_out_valid),
    .io_data_0_out_bits(PE_126_io_data_0_out_bits),
    .io_sig_stat2trans(PE_126_io_sig_stat2trans)
  );
  PE PE_127 ( // @[pearray.scala 101:13]
    .clock(PE_127_clock),
    .reset(PE_127_reset),
    .io_data_2_in_bits(PE_127_io_data_2_in_bits),
    .io_data_2_out_bits(PE_127_io_data_2_out_bits),
    .io_data_1_in_valid(PE_127_io_data_1_in_valid),
    .io_data_1_in_bits(PE_127_io_data_1_in_bits),
    .io_data_1_out_valid(PE_127_io_data_1_out_valid),
    .io_data_1_out_bits(PE_127_io_data_1_out_bits),
    .io_data_0_in_valid(PE_127_io_data_0_in_valid),
    .io_data_0_in_bits(PE_127_io_data_0_in_bits),
    .io_data_0_out_valid(PE_127_io_data_0_out_valid),
    .io_data_0_out_bits(PE_127_io_data_0_out_bits),
    .io_sig_stat2trans(PE_127_io_sig_stat2trans)
  );
  PENetwork PENetwork ( // @[pearray.scala 134:13]
    .io_to_pes_0_out_valid(PENetwork_io_to_pes_0_out_valid),
    .io_to_pes_0_out_bits(PENetwork_io_to_pes_0_out_bits),
    .io_to_pes_1_in_valid(PENetwork_io_to_pes_1_in_valid),
    .io_to_pes_1_in_bits(PENetwork_io_to_pes_1_in_bits),
    .io_to_pes_1_out_valid(PENetwork_io_to_pes_1_out_valid),
    .io_to_pes_1_out_bits(PENetwork_io_to_pes_1_out_bits),
    .io_to_pes_2_in_valid(PENetwork_io_to_pes_2_in_valid),
    .io_to_pes_2_in_bits(PENetwork_io_to_pes_2_in_bits),
    .io_to_pes_2_out_valid(PENetwork_io_to_pes_2_out_valid),
    .io_to_pes_2_out_bits(PENetwork_io_to_pes_2_out_bits),
    .io_to_pes_3_in_valid(PENetwork_io_to_pes_3_in_valid),
    .io_to_pes_3_in_bits(PENetwork_io_to_pes_3_in_bits),
    .io_to_pes_3_out_valid(PENetwork_io_to_pes_3_out_valid),
    .io_to_pes_3_out_bits(PENetwork_io_to_pes_3_out_bits),
    .io_to_pes_4_in_valid(PENetwork_io_to_pes_4_in_valid),
    .io_to_pes_4_in_bits(PENetwork_io_to_pes_4_in_bits),
    .io_to_pes_4_out_valid(PENetwork_io_to_pes_4_out_valid),
    .io_to_pes_4_out_bits(PENetwork_io_to_pes_4_out_bits),
    .io_to_pes_5_in_valid(PENetwork_io_to_pes_5_in_valid),
    .io_to_pes_5_in_bits(PENetwork_io_to_pes_5_in_bits),
    .io_to_pes_5_out_valid(PENetwork_io_to_pes_5_out_valid),
    .io_to_pes_5_out_bits(PENetwork_io_to_pes_5_out_bits),
    .io_to_pes_6_in_valid(PENetwork_io_to_pes_6_in_valid),
    .io_to_pes_6_in_bits(PENetwork_io_to_pes_6_in_bits),
    .io_to_pes_6_out_valid(PENetwork_io_to_pes_6_out_valid),
    .io_to_pes_6_out_bits(PENetwork_io_to_pes_6_out_bits),
    .io_to_pes_7_in_valid(PENetwork_io_to_pes_7_in_valid),
    .io_to_pes_7_in_bits(PENetwork_io_to_pes_7_in_bits),
    .io_to_pes_7_out_valid(PENetwork_io_to_pes_7_out_valid),
    .io_to_pes_7_out_bits(PENetwork_io_to_pes_7_out_bits),
    .io_to_mem_valid(PENetwork_io_to_mem_valid),
    .io_to_mem_bits(PENetwork_io_to_mem_bits)
  );
  PENetwork PENetwork_1 ( // @[pearray.scala 134:13]
    .io_to_pes_0_out_valid(PENetwork_1_io_to_pes_0_out_valid),
    .io_to_pes_0_out_bits(PENetwork_1_io_to_pes_0_out_bits),
    .io_to_pes_1_in_valid(PENetwork_1_io_to_pes_1_in_valid),
    .io_to_pes_1_in_bits(PENetwork_1_io_to_pes_1_in_bits),
    .io_to_pes_1_out_valid(PENetwork_1_io_to_pes_1_out_valid),
    .io_to_pes_1_out_bits(PENetwork_1_io_to_pes_1_out_bits),
    .io_to_pes_2_in_valid(PENetwork_1_io_to_pes_2_in_valid),
    .io_to_pes_2_in_bits(PENetwork_1_io_to_pes_2_in_bits),
    .io_to_pes_2_out_valid(PENetwork_1_io_to_pes_2_out_valid),
    .io_to_pes_2_out_bits(PENetwork_1_io_to_pes_2_out_bits),
    .io_to_pes_3_in_valid(PENetwork_1_io_to_pes_3_in_valid),
    .io_to_pes_3_in_bits(PENetwork_1_io_to_pes_3_in_bits),
    .io_to_pes_3_out_valid(PENetwork_1_io_to_pes_3_out_valid),
    .io_to_pes_3_out_bits(PENetwork_1_io_to_pes_3_out_bits),
    .io_to_pes_4_in_valid(PENetwork_1_io_to_pes_4_in_valid),
    .io_to_pes_4_in_bits(PENetwork_1_io_to_pes_4_in_bits),
    .io_to_pes_4_out_valid(PENetwork_1_io_to_pes_4_out_valid),
    .io_to_pes_4_out_bits(PENetwork_1_io_to_pes_4_out_bits),
    .io_to_pes_5_in_valid(PENetwork_1_io_to_pes_5_in_valid),
    .io_to_pes_5_in_bits(PENetwork_1_io_to_pes_5_in_bits),
    .io_to_pes_5_out_valid(PENetwork_1_io_to_pes_5_out_valid),
    .io_to_pes_5_out_bits(PENetwork_1_io_to_pes_5_out_bits),
    .io_to_pes_6_in_valid(PENetwork_1_io_to_pes_6_in_valid),
    .io_to_pes_6_in_bits(PENetwork_1_io_to_pes_6_in_bits),
    .io_to_pes_6_out_valid(PENetwork_1_io_to_pes_6_out_valid),
    .io_to_pes_6_out_bits(PENetwork_1_io_to_pes_6_out_bits),
    .io_to_pes_7_in_valid(PENetwork_1_io_to_pes_7_in_valid),
    .io_to_pes_7_in_bits(PENetwork_1_io_to_pes_7_in_bits),
    .io_to_pes_7_out_valid(PENetwork_1_io_to_pes_7_out_valid),
    .io_to_pes_7_out_bits(PENetwork_1_io_to_pes_7_out_bits),
    .io_to_mem_valid(PENetwork_1_io_to_mem_valid),
    .io_to_mem_bits(PENetwork_1_io_to_mem_bits)
  );
  PENetwork PENetwork_2 ( // @[pearray.scala 134:13]
    .io_to_pes_0_out_valid(PENetwork_2_io_to_pes_0_out_valid),
    .io_to_pes_0_out_bits(PENetwork_2_io_to_pes_0_out_bits),
    .io_to_pes_1_in_valid(PENetwork_2_io_to_pes_1_in_valid),
    .io_to_pes_1_in_bits(PENetwork_2_io_to_pes_1_in_bits),
    .io_to_pes_1_out_valid(PENetwork_2_io_to_pes_1_out_valid),
    .io_to_pes_1_out_bits(PENetwork_2_io_to_pes_1_out_bits),
    .io_to_pes_2_in_valid(PENetwork_2_io_to_pes_2_in_valid),
    .io_to_pes_2_in_bits(PENetwork_2_io_to_pes_2_in_bits),
    .io_to_pes_2_out_valid(PENetwork_2_io_to_pes_2_out_valid),
    .io_to_pes_2_out_bits(PENetwork_2_io_to_pes_2_out_bits),
    .io_to_pes_3_in_valid(PENetwork_2_io_to_pes_3_in_valid),
    .io_to_pes_3_in_bits(PENetwork_2_io_to_pes_3_in_bits),
    .io_to_pes_3_out_valid(PENetwork_2_io_to_pes_3_out_valid),
    .io_to_pes_3_out_bits(PENetwork_2_io_to_pes_3_out_bits),
    .io_to_pes_4_in_valid(PENetwork_2_io_to_pes_4_in_valid),
    .io_to_pes_4_in_bits(PENetwork_2_io_to_pes_4_in_bits),
    .io_to_pes_4_out_valid(PENetwork_2_io_to_pes_4_out_valid),
    .io_to_pes_4_out_bits(PENetwork_2_io_to_pes_4_out_bits),
    .io_to_pes_5_in_valid(PENetwork_2_io_to_pes_5_in_valid),
    .io_to_pes_5_in_bits(PENetwork_2_io_to_pes_5_in_bits),
    .io_to_pes_5_out_valid(PENetwork_2_io_to_pes_5_out_valid),
    .io_to_pes_5_out_bits(PENetwork_2_io_to_pes_5_out_bits),
    .io_to_pes_6_in_valid(PENetwork_2_io_to_pes_6_in_valid),
    .io_to_pes_6_in_bits(PENetwork_2_io_to_pes_6_in_bits),
    .io_to_pes_6_out_valid(PENetwork_2_io_to_pes_6_out_valid),
    .io_to_pes_6_out_bits(PENetwork_2_io_to_pes_6_out_bits),
    .io_to_pes_7_in_valid(PENetwork_2_io_to_pes_7_in_valid),
    .io_to_pes_7_in_bits(PENetwork_2_io_to_pes_7_in_bits),
    .io_to_pes_7_out_valid(PENetwork_2_io_to_pes_7_out_valid),
    .io_to_pes_7_out_bits(PENetwork_2_io_to_pes_7_out_bits),
    .io_to_mem_valid(PENetwork_2_io_to_mem_valid),
    .io_to_mem_bits(PENetwork_2_io_to_mem_bits)
  );
  PENetwork PENetwork_3 ( // @[pearray.scala 134:13]
    .io_to_pes_0_out_valid(PENetwork_3_io_to_pes_0_out_valid),
    .io_to_pes_0_out_bits(PENetwork_3_io_to_pes_0_out_bits),
    .io_to_pes_1_in_valid(PENetwork_3_io_to_pes_1_in_valid),
    .io_to_pes_1_in_bits(PENetwork_3_io_to_pes_1_in_bits),
    .io_to_pes_1_out_valid(PENetwork_3_io_to_pes_1_out_valid),
    .io_to_pes_1_out_bits(PENetwork_3_io_to_pes_1_out_bits),
    .io_to_pes_2_in_valid(PENetwork_3_io_to_pes_2_in_valid),
    .io_to_pes_2_in_bits(PENetwork_3_io_to_pes_2_in_bits),
    .io_to_pes_2_out_valid(PENetwork_3_io_to_pes_2_out_valid),
    .io_to_pes_2_out_bits(PENetwork_3_io_to_pes_2_out_bits),
    .io_to_pes_3_in_valid(PENetwork_3_io_to_pes_3_in_valid),
    .io_to_pes_3_in_bits(PENetwork_3_io_to_pes_3_in_bits),
    .io_to_pes_3_out_valid(PENetwork_3_io_to_pes_3_out_valid),
    .io_to_pes_3_out_bits(PENetwork_3_io_to_pes_3_out_bits),
    .io_to_pes_4_in_valid(PENetwork_3_io_to_pes_4_in_valid),
    .io_to_pes_4_in_bits(PENetwork_3_io_to_pes_4_in_bits),
    .io_to_pes_4_out_valid(PENetwork_3_io_to_pes_4_out_valid),
    .io_to_pes_4_out_bits(PENetwork_3_io_to_pes_4_out_bits),
    .io_to_pes_5_in_valid(PENetwork_3_io_to_pes_5_in_valid),
    .io_to_pes_5_in_bits(PENetwork_3_io_to_pes_5_in_bits),
    .io_to_pes_5_out_valid(PENetwork_3_io_to_pes_5_out_valid),
    .io_to_pes_5_out_bits(PENetwork_3_io_to_pes_5_out_bits),
    .io_to_pes_6_in_valid(PENetwork_3_io_to_pes_6_in_valid),
    .io_to_pes_6_in_bits(PENetwork_3_io_to_pes_6_in_bits),
    .io_to_pes_6_out_valid(PENetwork_3_io_to_pes_6_out_valid),
    .io_to_pes_6_out_bits(PENetwork_3_io_to_pes_6_out_bits),
    .io_to_pes_7_in_valid(PENetwork_3_io_to_pes_7_in_valid),
    .io_to_pes_7_in_bits(PENetwork_3_io_to_pes_7_in_bits),
    .io_to_pes_7_out_valid(PENetwork_3_io_to_pes_7_out_valid),
    .io_to_pes_7_out_bits(PENetwork_3_io_to_pes_7_out_bits),
    .io_to_mem_valid(PENetwork_3_io_to_mem_valid),
    .io_to_mem_bits(PENetwork_3_io_to_mem_bits)
  );
  PENetwork PENetwork_4 ( // @[pearray.scala 134:13]
    .io_to_pes_0_out_valid(PENetwork_4_io_to_pes_0_out_valid),
    .io_to_pes_0_out_bits(PENetwork_4_io_to_pes_0_out_bits),
    .io_to_pes_1_in_valid(PENetwork_4_io_to_pes_1_in_valid),
    .io_to_pes_1_in_bits(PENetwork_4_io_to_pes_1_in_bits),
    .io_to_pes_1_out_valid(PENetwork_4_io_to_pes_1_out_valid),
    .io_to_pes_1_out_bits(PENetwork_4_io_to_pes_1_out_bits),
    .io_to_pes_2_in_valid(PENetwork_4_io_to_pes_2_in_valid),
    .io_to_pes_2_in_bits(PENetwork_4_io_to_pes_2_in_bits),
    .io_to_pes_2_out_valid(PENetwork_4_io_to_pes_2_out_valid),
    .io_to_pes_2_out_bits(PENetwork_4_io_to_pes_2_out_bits),
    .io_to_pes_3_in_valid(PENetwork_4_io_to_pes_3_in_valid),
    .io_to_pes_3_in_bits(PENetwork_4_io_to_pes_3_in_bits),
    .io_to_pes_3_out_valid(PENetwork_4_io_to_pes_3_out_valid),
    .io_to_pes_3_out_bits(PENetwork_4_io_to_pes_3_out_bits),
    .io_to_pes_4_in_valid(PENetwork_4_io_to_pes_4_in_valid),
    .io_to_pes_4_in_bits(PENetwork_4_io_to_pes_4_in_bits),
    .io_to_pes_4_out_valid(PENetwork_4_io_to_pes_4_out_valid),
    .io_to_pes_4_out_bits(PENetwork_4_io_to_pes_4_out_bits),
    .io_to_pes_5_in_valid(PENetwork_4_io_to_pes_5_in_valid),
    .io_to_pes_5_in_bits(PENetwork_4_io_to_pes_5_in_bits),
    .io_to_pes_5_out_valid(PENetwork_4_io_to_pes_5_out_valid),
    .io_to_pes_5_out_bits(PENetwork_4_io_to_pes_5_out_bits),
    .io_to_pes_6_in_valid(PENetwork_4_io_to_pes_6_in_valid),
    .io_to_pes_6_in_bits(PENetwork_4_io_to_pes_6_in_bits),
    .io_to_pes_6_out_valid(PENetwork_4_io_to_pes_6_out_valid),
    .io_to_pes_6_out_bits(PENetwork_4_io_to_pes_6_out_bits),
    .io_to_pes_7_in_valid(PENetwork_4_io_to_pes_7_in_valid),
    .io_to_pes_7_in_bits(PENetwork_4_io_to_pes_7_in_bits),
    .io_to_pes_7_out_valid(PENetwork_4_io_to_pes_7_out_valid),
    .io_to_pes_7_out_bits(PENetwork_4_io_to_pes_7_out_bits),
    .io_to_mem_valid(PENetwork_4_io_to_mem_valid),
    .io_to_mem_bits(PENetwork_4_io_to_mem_bits)
  );
  PENetwork PENetwork_5 ( // @[pearray.scala 134:13]
    .io_to_pes_0_out_valid(PENetwork_5_io_to_pes_0_out_valid),
    .io_to_pes_0_out_bits(PENetwork_5_io_to_pes_0_out_bits),
    .io_to_pes_1_in_valid(PENetwork_5_io_to_pes_1_in_valid),
    .io_to_pes_1_in_bits(PENetwork_5_io_to_pes_1_in_bits),
    .io_to_pes_1_out_valid(PENetwork_5_io_to_pes_1_out_valid),
    .io_to_pes_1_out_bits(PENetwork_5_io_to_pes_1_out_bits),
    .io_to_pes_2_in_valid(PENetwork_5_io_to_pes_2_in_valid),
    .io_to_pes_2_in_bits(PENetwork_5_io_to_pes_2_in_bits),
    .io_to_pes_2_out_valid(PENetwork_5_io_to_pes_2_out_valid),
    .io_to_pes_2_out_bits(PENetwork_5_io_to_pes_2_out_bits),
    .io_to_pes_3_in_valid(PENetwork_5_io_to_pes_3_in_valid),
    .io_to_pes_3_in_bits(PENetwork_5_io_to_pes_3_in_bits),
    .io_to_pes_3_out_valid(PENetwork_5_io_to_pes_3_out_valid),
    .io_to_pes_3_out_bits(PENetwork_5_io_to_pes_3_out_bits),
    .io_to_pes_4_in_valid(PENetwork_5_io_to_pes_4_in_valid),
    .io_to_pes_4_in_bits(PENetwork_5_io_to_pes_4_in_bits),
    .io_to_pes_4_out_valid(PENetwork_5_io_to_pes_4_out_valid),
    .io_to_pes_4_out_bits(PENetwork_5_io_to_pes_4_out_bits),
    .io_to_pes_5_in_valid(PENetwork_5_io_to_pes_5_in_valid),
    .io_to_pes_5_in_bits(PENetwork_5_io_to_pes_5_in_bits),
    .io_to_pes_5_out_valid(PENetwork_5_io_to_pes_5_out_valid),
    .io_to_pes_5_out_bits(PENetwork_5_io_to_pes_5_out_bits),
    .io_to_pes_6_in_valid(PENetwork_5_io_to_pes_6_in_valid),
    .io_to_pes_6_in_bits(PENetwork_5_io_to_pes_6_in_bits),
    .io_to_pes_6_out_valid(PENetwork_5_io_to_pes_6_out_valid),
    .io_to_pes_6_out_bits(PENetwork_5_io_to_pes_6_out_bits),
    .io_to_pes_7_in_valid(PENetwork_5_io_to_pes_7_in_valid),
    .io_to_pes_7_in_bits(PENetwork_5_io_to_pes_7_in_bits),
    .io_to_pes_7_out_valid(PENetwork_5_io_to_pes_7_out_valid),
    .io_to_pes_7_out_bits(PENetwork_5_io_to_pes_7_out_bits),
    .io_to_mem_valid(PENetwork_5_io_to_mem_valid),
    .io_to_mem_bits(PENetwork_5_io_to_mem_bits)
  );
  PENetwork PENetwork_6 ( // @[pearray.scala 134:13]
    .io_to_pes_0_out_valid(PENetwork_6_io_to_pes_0_out_valid),
    .io_to_pes_0_out_bits(PENetwork_6_io_to_pes_0_out_bits),
    .io_to_pes_1_in_valid(PENetwork_6_io_to_pes_1_in_valid),
    .io_to_pes_1_in_bits(PENetwork_6_io_to_pes_1_in_bits),
    .io_to_pes_1_out_valid(PENetwork_6_io_to_pes_1_out_valid),
    .io_to_pes_1_out_bits(PENetwork_6_io_to_pes_1_out_bits),
    .io_to_pes_2_in_valid(PENetwork_6_io_to_pes_2_in_valid),
    .io_to_pes_2_in_bits(PENetwork_6_io_to_pes_2_in_bits),
    .io_to_pes_2_out_valid(PENetwork_6_io_to_pes_2_out_valid),
    .io_to_pes_2_out_bits(PENetwork_6_io_to_pes_2_out_bits),
    .io_to_pes_3_in_valid(PENetwork_6_io_to_pes_3_in_valid),
    .io_to_pes_3_in_bits(PENetwork_6_io_to_pes_3_in_bits),
    .io_to_pes_3_out_valid(PENetwork_6_io_to_pes_3_out_valid),
    .io_to_pes_3_out_bits(PENetwork_6_io_to_pes_3_out_bits),
    .io_to_pes_4_in_valid(PENetwork_6_io_to_pes_4_in_valid),
    .io_to_pes_4_in_bits(PENetwork_6_io_to_pes_4_in_bits),
    .io_to_pes_4_out_valid(PENetwork_6_io_to_pes_4_out_valid),
    .io_to_pes_4_out_bits(PENetwork_6_io_to_pes_4_out_bits),
    .io_to_pes_5_in_valid(PENetwork_6_io_to_pes_5_in_valid),
    .io_to_pes_5_in_bits(PENetwork_6_io_to_pes_5_in_bits),
    .io_to_pes_5_out_valid(PENetwork_6_io_to_pes_5_out_valid),
    .io_to_pes_5_out_bits(PENetwork_6_io_to_pes_5_out_bits),
    .io_to_pes_6_in_valid(PENetwork_6_io_to_pes_6_in_valid),
    .io_to_pes_6_in_bits(PENetwork_6_io_to_pes_6_in_bits),
    .io_to_pes_6_out_valid(PENetwork_6_io_to_pes_6_out_valid),
    .io_to_pes_6_out_bits(PENetwork_6_io_to_pes_6_out_bits),
    .io_to_pes_7_in_valid(PENetwork_6_io_to_pes_7_in_valid),
    .io_to_pes_7_in_bits(PENetwork_6_io_to_pes_7_in_bits),
    .io_to_pes_7_out_valid(PENetwork_6_io_to_pes_7_out_valid),
    .io_to_pes_7_out_bits(PENetwork_6_io_to_pes_7_out_bits),
    .io_to_mem_valid(PENetwork_6_io_to_mem_valid),
    .io_to_mem_bits(PENetwork_6_io_to_mem_bits)
  );
  PENetwork PENetwork_7 ( // @[pearray.scala 134:13]
    .io_to_pes_0_out_valid(PENetwork_7_io_to_pes_0_out_valid),
    .io_to_pes_0_out_bits(PENetwork_7_io_to_pes_0_out_bits),
    .io_to_pes_1_in_valid(PENetwork_7_io_to_pes_1_in_valid),
    .io_to_pes_1_in_bits(PENetwork_7_io_to_pes_1_in_bits),
    .io_to_pes_1_out_valid(PENetwork_7_io_to_pes_1_out_valid),
    .io_to_pes_1_out_bits(PENetwork_7_io_to_pes_1_out_bits),
    .io_to_pes_2_in_valid(PENetwork_7_io_to_pes_2_in_valid),
    .io_to_pes_2_in_bits(PENetwork_7_io_to_pes_2_in_bits),
    .io_to_pes_2_out_valid(PENetwork_7_io_to_pes_2_out_valid),
    .io_to_pes_2_out_bits(PENetwork_7_io_to_pes_2_out_bits),
    .io_to_pes_3_in_valid(PENetwork_7_io_to_pes_3_in_valid),
    .io_to_pes_3_in_bits(PENetwork_7_io_to_pes_3_in_bits),
    .io_to_pes_3_out_valid(PENetwork_7_io_to_pes_3_out_valid),
    .io_to_pes_3_out_bits(PENetwork_7_io_to_pes_3_out_bits),
    .io_to_pes_4_in_valid(PENetwork_7_io_to_pes_4_in_valid),
    .io_to_pes_4_in_bits(PENetwork_7_io_to_pes_4_in_bits),
    .io_to_pes_4_out_valid(PENetwork_7_io_to_pes_4_out_valid),
    .io_to_pes_4_out_bits(PENetwork_7_io_to_pes_4_out_bits),
    .io_to_pes_5_in_valid(PENetwork_7_io_to_pes_5_in_valid),
    .io_to_pes_5_in_bits(PENetwork_7_io_to_pes_5_in_bits),
    .io_to_pes_5_out_valid(PENetwork_7_io_to_pes_5_out_valid),
    .io_to_pes_5_out_bits(PENetwork_7_io_to_pes_5_out_bits),
    .io_to_pes_6_in_valid(PENetwork_7_io_to_pes_6_in_valid),
    .io_to_pes_6_in_bits(PENetwork_7_io_to_pes_6_in_bits),
    .io_to_pes_6_out_valid(PENetwork_7_io_to_pes_6_out_valid),
    .io_to_pes_6_out_bits(PENetwork_7_io_to_pes_6_out_bits),
    .io_to_pes_7_in_valid(PENetwork_7_io_to_pes_7_in_valid),
    .io_to_pes_7_in_bits(PENetwork_7_io_to_pes_7_in_bits),
    .io_to_pes_7_out_valid(PENetwork_7_io_to_pes_7_out_valid),
    .io_to_pes_7_out_bits(PENetwork_7_io_to_pes_7_out_bits),
    .io_to_mem_valid(PENetwork_7_io_to_mem_valid),
    .io_to_mem_bits(PENetwork_7_io_to_mem_bits)
  );
  PENetwork PENetwork_8 ( // @[pearray.scala 134:13]
    .io_to_pes_0_out_valid(PENetwork_8_io_to_pes_0_out_valid),
    .io_to_pes_0_out_bits(PENetwork_8_io_to_pes_0_out_bits),
    .io_to_pes_1_in_valid(PENetwork_8_io_to_pes_1_in_valid),
    .io_to_pes_1_in_bits(PENetwork_8_io_to_pes_1_in_bits),
    .io_to_pes_1_out_valid(PENetwork_8_io_to_pes_1_out_valid),
    .io_to_pes_1_out_bits(PENetwork_8_io_to_pes_1_out_bits),
    .io_to_pes_2_in_valid(PENetwork_8_io_to_pes_2_in_valid),
    .io_to_pes_2_in_bits(PENetwork_8_io_to_pes_2_in_bits),
    .io_to_pes_2_out_valid(PENetwork_8_io_to_pes_2_out_valid),
    .io_to_pes_2_out_bits(PENetwork_8_io_to_pes_2_out_bits),
    .io_to_pes_3_in_valid(PENetwork_8_io_to_pes_3_in_valid),
    .io_to_pes_3_in_bits(PENetwork_8_io_to_pes_3_in_bits),
    .io_to_pes_3_out_valid(PENetwork_8_io_to_pes_3_out_valid),
    .io_to_pes_3_out_bits(PENetwork_8_io_to_pes_3_out_bits),
    .io_to_pes_4_in_valid(PENetwork_8_io_to_pes_4_in_valid),
    .io_to_pes_4_in_bits(PENetwork_8_io_to_pes_4_in_bits),
    .io_to_pes_4_out_valid(PENetwork_8_io_to_pes_4_out_valid),
    .io_to_pes_4_out_bits(PENetwork_8_io_to_pes_4_out_bits),
    .io_to_pes_5_in_valid(PENetwork_8_io_to_pes_5_in_valid),
    .io_to_pes_5_in_bits(PENetwork_8_io_to_pes_5_in_bits),
    .io_to_pes_5_out_valid(PENetwork_8_io_to_pes_5_out_valid),
    .io_to_pes_5_out_bits(PENetwork_8_io_to_pes_5_out_bits),
    .io_to_pes_6_in_valid(PENetwork_8_io_to_pes_6_in_valid),
    .io_to_pes_6_in_bits(PENetwork_8_io_to_pes_6_in_bits),
    .io_to_pes_6_out_valid(PENetwork_8_io_to_pes_6_out_valid),
    .io_to_pes_6_out_bits(PENetwork_8_io_to_pes_6_out_bits),
    .io_to_pes_7_in_valid(PENetwork_8_io_to_pes_7_in_valid),
    .io_to_pes_7_in_bits(PENetwork_8_io_to_pes_7_in_bits),
    .io_to_pes_7_out_valid(PENetwork_8_io_to_pes_7_out_valid),
    .io_to_pes_7_out_bits(PENetwork_8_io_to_pes_7_out_bits),
    .io_to_mem_valid(PENetwork_8_io_to_mem_valid),
    .io_to_mem_bits(PENetwork_8_io_to_mem_bits)
  );
  PENetwork PENetwork_9 ( // @[pearray.scala 134:13]
    .io_to_pes_0_out_valid(PENetwork_9_io_to_pes_0_out_valid),
    .io_to_pes_0_out_bits(PENetwork_9_io_to_pes_0_out_bits),
    .io_to_pes_1_in_valid(PENetwork_9_io_to_pes_1_in_valid),
    .io_to_pes_1_in_bits(PENetwork_9_io_to_pes_1_in_bits),
    .io_to_pes_1_out_valid(PENetwork_9_io_to_pes_1_out_valid),
    .io_to_pes_1_out_bits(PENetwork_9_io_to_pes_1_out_bits),
    .io_to_pes_2_in_valid(PENetwork_9_io_to_pes_2_in_valid),
    .io_to_pes_2_in_bits(PENetwork_9_io_to_pes_2_in_bits),
    .io_to_pes_2_out_valid(PENetwork_9_io_to_pes_2_out_valid),
    .io_to_pes_2_out_bits(PENetwork_9_io_to_pes_2_out_bits),
    .io_to_pes_3_in_valid(PENetwork_9_io_to_pes_3_in_valid),
    .io_to_pes_3_in_bits(PENetwork_9_io_to_pes_3_in_bits),
    .io_to_pes_3_out_valid(PENetwork_9_io_to_pes_3_out_valid),
    .io_to_pes_3_out_bits(PENetwork_9_io_to_pes_3_out_bits),
    .io_to_pes_4_in_valid(PENetwork_9_io_to_pes_4_in_valid),
    .io_to_pes_4_in_bits(PENetwork_9_io_to_pes_4_in_bits),
    .io_to_pes_4_out_valid(PENetwork_9_io_to_pes_4_out_valid),
    .io_to_pes_4_out_bits(PENetwork_9_io_to_pes_4_out_bits),
    .io_to_pes_5_in_valid(PENetwork_9_io_to_pes_5_in_valid),
    .io_to_pes_5_in_bits(PENetwork_9_io_to_pes_5_in_bits),
    .io_to_pes_5_out_valid(PENetwork_9_io_to_pes_5_out_valid),
    .io_to_pes_5_out_bits(PENetwork_9_io_to_pes_5_out_bits),
    .io_to_pes_6_in_valid(PENetwork_9_io_to_pes_6_in_valid),
    .io_to_pes_6_in_bits(PENetwork_9_io_to_pes_6_in_bits),
    .io_to_pes_6_out_valid(PENetwork_9_io_to_pes_6_out_valid),
    .io_to_pes_6_out_bits(PENetwork_9_io_to_pes_6_out_bits),
    .io_to_pes_7_in_valid(PENetwork_9_io_to_pes_7_in_valid),
    .io_to_pes_7_in_bits(PENetwork_9_io_to_pes_7_in_bits),
    .io_to_pes_7_out_valid(PENetwork_9_io_to_pes_7_out_valid),
    .io_to_pes_7_out_bits(PENetwork_9_io_to_pes_7_out_bits),
    .io_to_mem_valid(PENetwork_9_io_to_mem_valid),
    .io_to_mem_bits(PENetwork_9_io_to_mem_bits)
  );
  PENetwork PENetwork_10 ( // @[pearray.scala 134:13]
    .io_to_pes_0_out_valid(PENetwork_10_io_to_pes_0_out_valid),
    .io_to_pes_0_out_bits(PENetwork_10_io_to_pes_0_out_bits),
    .io_to_pes_1_in_valid(PENetwork_10_io_to_pes_1_in_valid),
    .io_to_pes_1_in_bits(PENetwork_10_io_to_pes_1_in_bits),
    .io_to_pes_1_out_valid(PENetwork_10_io_to_pes_1_out_valid),
    .io_to_pes_1_out_bits(PENetwork_10_io_to_pes_1_out_bits),
    .io_to_pes_2_in_valid(PENetwork_10_io_to_pes_2_in_valid),
    .io_to_pes_2_in_bits(PENetwork_10_io_to_pes_2_in_bits),
    .io_to_pes_2_out_valid(PENetwork_10_io_to_pes_2_out_valid),
    .io_to_pes_2_out_bits(PENetwork_10_io_to_pes_2_out_bits),
    .io_to_pes_3_in_valid(PENetwork_10_io_to_pes_3_in_valid),
    .io_to_pes_3_in_bits(PENetwork_10_io_to_pes_3_in_bits),
    .io_to_pes_3_out_valid(PENetwork_10_io_to_pes_3_out_valid),
    .io_to_pes_3_out_bits(PENetwork_10_io_to_pes_3_out_bits),
    .io_to_pes_4_in_valid(PENetwork_10_io_to_pes_4_in_valid),
    .io_to_pes_4_in_bits(PENetwork_10_io_to_pes_4_in_bits),
    .io_to_pes_4_out_valid(PENetwork_10_io_to_pes_4_out_valid),
    .io_to_pes_4_out_bits(PENetwork_10_io_to_pes_4_out_bits),
    .io_to_pes_5_in_valid(PENetwork_10_io_to_pes_5_in_valid),
    .io_to_pes_5_in_bits(PENetwork_10_io_to_pes_5_in_bits),
    .io_to_pes_5_out_valid(PENetwork_10_io_to_pes_5_out_valid),
    .io_to_pes_5_out_bits(PENetwork_10_io_to_pes_5_out_bits),
    .io_to_pes_6_in_valid(PENetwork_10_io_to_pes_6_in_valid),
    .io_to_pes_6_in_bits(PENetwork_10_io_to_pes_6_in_bits),
    .io_to_pes_6_out_valid(PENetwork_10_io_to_pes_6_out_valid),
    .io_to_pes_6_out_bits(PENetwork_10_io_to_pes_6_out_bits),
    .io_to_pes_7_in_valid(PENetwork_10_io_to_pes_7_in_valid),
    .io_to_pes_7_in_bits(PENetwork_10_io_to_pes_7_in_bits),
    .io_to_pes_7_out_valid(PENetwork_10_io_to_pes_7_out_valid),
    .io_to_pes_7_out_bits(PENetwork_10_io_to_pes_7_out_bits),
    .io_to_mem_valid(PENetwork_10_io_to_mem_valid),
    .io_to_mem_bits(PENetwork_10_io_to_mem_bits)
  );
  PENetwork PENetwork_11 ( // @[pearray.scala 134:13]
    .io_to_pes_0_out_valid(PENetwork_11_io_to_pes_0_out_valid),
    .io_to_pes_0_out_bits(PENetwork_11_io_to_pes_0_out_bits),
    .io_to_pes_1_in_valid(PENetwork_11_io_to_pes_1_in_valid),
    .io_to_pes_1_in_bits(PENetwork_11_io_to_pes_1_in_bits),
    .io_to_pes_1_out_valid(PENetwork_11_io_to_pes_1_out_valid),
    .io_to_pes_1_out_bits(PENetwork_11_io_to_pes_1_out_bits),
    .io_to_pes_2_in_valid(PENetwork_11_io_to_pes_2_in_valid),
    .io_to_pes_2_in_bits(PENetwork_11_io_to_pes_2_in_bits),
    .io_to_pes_2_out_valid(PENetwork_11_io_to_pes_2_out_valid),
    .io_to_pes_2_out_bits(PENetwork_11_io_to_pes_2_out_bits),
    .io_to_pes_3_in_valid(PENetwork_11_io_to_pes_3_in_valid),
    .io_to_pes_3_in_bits(PENetwork_11_io_to_pes_3_in_bits),
    .io_to_pes_3_out_valid(PENetwork_11_io_to_pes_3_out_valid),
    .io_to_pes_3_out_bits(PENetwork_11_io_to_pes_3_out_bits),
    .io_to_pes_4_in_valid(PENetwork_11_io_to_pes_4_in_valid),
    .io_to_pes_4_in_bits(PENetwork_11_io_to_pes_4_in_bits),
    .io_to_pes_4_out_valid(PENetwork_11_io_to_pes_4_out_valid),
    .io_to_pes_4_out_bits(PENetwork_11_io_to_pes_4_out_bits),
    .io_to_pes_5_in_valid(PENetwork_11_io_to_pes_5_in_valid),
    .io_to_pes_5_in_bits(PENetwork_11_io_to_pes_5_in_bits),
    .io_to_pes_5_out_valid(PENetwork_11_io_to_pes_5_out_valid),
    .io_to_pes_5_out_bits(PENetwork_11_io_to_pes_5_out_bits),
    .io_to_pes_6_in_valid(PENetwork_11_io_to_pes_6_in_valid),
    .io_to_pes_6_in_bits(PENetwork_11_io_to_pes_6_in_bits),
    .io_to_pes_6_out_valid(PENetwork_11_io_to_pes_6_out_valid),
    .io_to_pes_6_out_bits(PENetwork_11_io_to_pes_6_out_bits),
    .io_to_pes_7_in_valid(PENetwork_11_io_to_pes_7_in_valid),
    .io_to_pes_7_in_bits(PENetwork_11_io_to_pes_7_in_bits),
    .io_to_pes_7_out_valid(PENetwork_11_io_to_pes_7_out_valid),
    .io_to_pes_7_out_bits(PENetwork_11_io_to_pes_7_out_bits),
    .io_to_mem_valid(PENetwork_11_io_to_mem_valid),
    .io_to_mem_bits(PENetwork_11_io_to_mem_bits)
  );
  PENetwork PENetwork_12 ( // @[pearray.scala 134:13]
    .io_to_pes_0_out_valid(PENetwork_12_io_to_pes_0_out_valid),
    .io_to_pes_0_out_bits(PENetwork_12_io_to_pes_0_out_bits),
    .io_to_pes_1_in_valid(PENetwork_12_io_to_pes_1_in_valid),
    .io_to_pes_1_in_bits(PENetwork_12_io_to_pes_1_in_bits),
    .io_to_pes_1_out_valid(PENetwork_12_io_to_pes_1_out_valid),
    .io_to_pes_1_out_bits(PENetwork_12_io_to_pes_1_out_bits),
    .io_to_pes_2_in_valid(PENetwork_12_io_to_pes_2_in_valid),
    .io_to_pes_2_in_bits(PENetwork_12_io_to_pes_2_in_bits),
    .io_to_pes_2_out_valid(PENetwork_12_io_to_pes_2_out_valid),
    .io_to_pes_2_out_bits(PENetwork_12_io_to_pes_2_out_bits),
    .io_to_pes_3_in_valid(PENetwork_12_io_to_pes_3_in_valid),
    .io_to_pes_3_in_bits(PENetwork_12_io_to_pes_3_in_bits),
    .io_to_pes_3_out_valid(PENetwork_12_io_to_pes_3_out_valid),
    .io_to_pes_3_out_bits(PENetwork_12_io_to_pes_3_out_bits),
    .io_to_pes_4_in_valid(PENetwork_12_io_to_pes_4_in_valid),
    .io_to_pes_4_in_bits(PENetwork_12_io_to_pes_4_in_bits),
    .io_to_pes_4_out_valid(PENetwork_12_io_to_pes_4_out_valid),
    .io_to_pes_4_out_bits(PENetwork_12_io_to_pes_4_out_bits),
    .io_to_pes_5_in_valid(PENetwork_12_io_to_pes_5_in_valid),
    .io_to_pes_5_in_bits(PENetwork_12_io_to_pes_5_in_bits),
    .io_to_pes_5_out_valid(PENetwork_12_io_to_pes_5_out_valid),
    .io_to_pes_5_out_bits(PENetwork_12_io_to_pes_5_out_bits),
    .io_to_pes_6_in_valid(PENetwork_12_io_to_pes_6_in_valid),
    .io_to_pes_6_in_bits(PENetwork_12_io_to_pes_6_in_bits),
    .io_to_pes_6_out_valid(PENetwork_12_io_to_pes_6_out_valid),
    .io_to_pes_6_out_bits(PENetwork_12_io_to_pes_6_out_bits),
    .io_to_pes_7_in_valid(PENetwork_12_io_to_pes_7_in_valid),
    .io_to_pes_7_in_bits(PENetwork_12_io_to_pes_7_in_bits),
    .io_to_pes_7_out_valid(PENetwork_12_io_to_pes_7_out_valid),
    .io_to_pes_7_out_bits(PENetwork_12_io_to_pes_7_out_bits),
    .io_to_mem_valid(PENetwork_12_io_to_mem_valid),
    .io_to_mem_bits(PENetwork_12_io_to_mem_bits)
  );
  PENetwork PENetwork_13 ( // @[pearray.scala 134:13]
    .io_to_pes_0_out_valid(PENetwork_13_io_to_pes_0_out_valid),
    .io_to_pes_0_out_bits(PENetwork_13_io_to_pes_0_out_bits),
    .io_to_pes_1_in_valid(PENetwork_13_io_to_pes_1_in_valid),
    .io_to_pes_1_in_bits(PENetwork_13_io_to_pes_1_in_bits),
    .io_to_pes_1_out_valid(PENetwork_13_io_to_pes_1_out_valid),
    .io_to_pes_1_out_bits(PENetwork_13_io_to_pes_1_out_bits),
    .io_to_pes_2_in_valid(PENetwork_13_io_to_pes_2_in_valid),
    .io_to_pes_2_in_bits(PENetwork_13_io_to_pes_2_in_bits),
    .io_to_pes_2_out_valid(PENetwork_13_io_to_pes_2_out_valid),
    .io_to_pes_2_out_bits(PENetwork_13_io_to_pes_2_out_bits),
    .io_to_pes_3_in_valid(PENetwork_13_io_to_pes_3_in_valid),
    .io_to_pes_3_in_bits(PENetwork_13_io_to_pes_3_in_bits),
    .io_to_pes_3_out_valid(PENetwork_13_io_to_pes_3_out_valid),
    .io_to_pes_3_out_bits(PENetwork_13_io_to_pes_3_out_bits),
    .io_to_pes_4_in_valid(PENetwork_13_io_to_pes_4_in_valid),
    .io_to_pes_4_in_bits(PENetwork_13_io_to_pes_4_in_bits),
    .io_to_pes_4_out_valid(PENetwork_13_io_to_pes_4_out_valid),
    .io_to_pes_4_out_bits(PENetwork_13_io_to_pes_4_out_bits),
    .io_to_pes_5_in_valid(PENetwork_13_io_to_pes_5_in_valid),
    .io_to_pes_5_in_bits(PENetwork_13_io_to_pes_5_in_bits),
    .io_to_pes_5_out_valid(PENetwork_13_io_to_pes_5_out_valid),
    .io_to_pes_5_out_bits(PENetwork_13_io_to_pes_5_out_bits),
    .io_to_pes_6_in_valid(PENetwork_13_io_to_pes_6_in_valid),
    .io_to_pes_6_in_bits(PENetwork_13_io_to_pes_6_in_bits),
    .io_to_pes_6_out_valid(PENetwork_13_io_to_pes_6_out_valid),
    .io_to_pes_6_out_bits(PENetwork_13_io_to_pes_6_out_bits),
    .io_to_pes_7_in_valid(PENetwork_13_io_to_pes_7_in_valid),
    .io_to_pes_7_in_bits(PENetwork_13_io_to_pes_7_in_bits),
    .io_to_pes_7_out_valid(PENetwork_13_io_to_pes_7_out_valid),
    .io_to_pes_7_out_bits(PENetwork_13_io_to_pes_7_out_bits),
    .io_to_mem_valid(PENetwork_13_io_to_mem_valid),
    .io_to_mem_bits(PENetwork_13_io_to_mem_bits)
  );
  PENetwork PENetwork_14 ( // @[pearray.scala 134:13]
    .io_to_pes_0_out_valid(PENetwork_14_io_to_pes_0_out_valid),
    .io_to_pes_0_out_bits(PENetwork_14_io_to_pes_0_out_bits),
    .io_to_pes_1_in_valid(PENetwork_14_io_to_pes_1_in_valid),
    .io_to_pes_1_in_bits(PENetwork_14_io_to_pes_1_in_bits),
    .io_to_pes_1_out_valid(PENetwork_14_io_to_pes_1_out_valid),
    .io_to_pes_1_out_bits(PENetwork_14_io_to_pes_1_out_bits),
    .io_to_pes_2_in_valid(PENetwork_14_io_to_pes_2_in_valid),
    .io_to_pes_2_in_bits(PENetwork_14_io_to_pes_2_in_bits),
    .io_to_pes_2_out_valid(PENetwork_14_io_to_pes_2_out_valid),
    .io_to_pes_2_out_bits(PENetwork_14_io_to_pes_2_out_bits),
    .io_to_pes_3_in_valid(PENetwork_14_io_to_pes_3_in_valid),
    .io_to_pes_3_in_bits(PENetwork_14_io_to_pes_3_in_bits),
    .io_to_pes_3_out_valid(PENetwork_14_io_to_pes_3_out_valid),
    .io_to_pes_3_out_bits(PENetwork_14_io_to_pes_3_out_bits),
    .io_to_pes_4_in_valid(PENetwork_14_io_to_pes_4_in_valid),
    .io_to_pes_4_in_bits(PENetwork_14_io_to_pes_4_in_bits),
    .io_to_pes_4_out_valid(PENetwork_14_io_to_pes_4_out_valid),
    .io_to_pes_4_out_bits(PENetwork_14_io_to_pes_4_out_bits),
    .io_to_pes_5_in_valid(PENetwork_14_io_to_pes_5_in_valid),
    .io_to_pes_5_in_bits(PENetwork_14_io_to_pes_5_in_bits),
    .io_to_pes_5_out_valid(PENetwork_14_io_to_pes_5_out_valid),
    .io_to_pes_5_out_bits(PENetwork_14_io_to_pes_5_out_bits),
    .io_to_pes_6_in_valid(PENetwork_14_io_to_pes_6_in_valid),
    .io_to_pes_6_in_bits(PENetwork_14_io_to_pes_6_in_bits),
    .io_to_pes_6_out_valid(PENetwork_14_io_to_pes_6_out_valid),
    .io_to_pes_6_out_bits(PENetwork_14_io_to_pes_6_out_bits),
    .io_to_pes_7_in_valid(PENetwork_14_io_to_pes_7_in_valid),
    .io_to_pes_7_in_bits(PENetwork_14_io_to_pes_7_in_bits),
    .io_to_pes_7_out_valid(PENetwork_14_io_to_pes_7_out_valid),
    .io_to_pes_7_out_bits(PENetwork_14_io_to_pes_7_out_bits),
    .io_to_mem_valid(PENetwork_14_io_to_mem_valid),
    .io_to_mem_bits(PENetwork_14_io_to_mem_bits)
  );
  PENetwork PENetwork_15 ( // @[pearray.scala 134:13]
    .io_to_pes_0_out_valid(PENetwork_15_io_to_pes_0_out_valid),
    .io_to_pes_0_out_bits(PENetwork_15_io_to_pes_0_out_bits),
    .io_to_pes_1_in_valid(PENetwork_15_io_to_pes_1_in_valid),
    .io_to_pes_1_in_bits(PENetwork_15_io_to_pes_1_in_bits),
    .io_to_pes_1_out_valid(PENetwork_15_io_to_pes_1_out_valid),
    .io_to_pes_1_out_bits(PENetwork_15_io_to_pes_1_out_bits),
    .io_to_pes_2_in_valid(PENetwork_15_io_to_pes_2_in_valid),
    .io_to_pes_2_in_bits(PENetwork_15_io_to_pes_2_in_bits),
    .io_to_pes_2_out_valid(PENetwork_15_io_to_pes_2_out_valid),
    .io_to_pes_2_out_bits(PENetwork_15_io_to_pes_2_out_bits),
    .io_to_pes_3_in_valid(PENetwork_15_io_to_pes_3_in_valid),
    .io_to_pes_3_in_bits(PENetwork_15_io_to_pes_3_in_bits),
    .io_to_pes_3_out_valid(PENetwork_15_io_to_pes_3_out_valid),
    .io_to_pes_3_out_bits(PENetwork_15_io_to_pes_3_out_bits),
    .io_to_pes_4_in_valid(PENetwork_15_io_to_pes_4_in_valid),
    .io_to_pes_4_in_bits(PENetwork_15_io_to_pes_4_in_bits),
    .io_to_pes_4_out_valid(PENetwork_15_io_to_pes_4_out_valid),
    .io_to_pes_4_out_bits(PENetwork_15_io_to_pes_4_out_bits),
    .io_to_pes_5_in_valid(PENetwork_15_io_to_pes_5_in_valid),
    .io_to_pes_5_in_bits(PENetwork_15_io_to_pes_5_in_bits),
    .io_to_pes_5_out_valid(PENetwork_15_io_to_pes_5_out_valid),
    .io_to_pes_5_out_bits(PENetwork_15_io_to_pes_5_out_bits),
    .io_to_pes_6_in_valid(PENetwork_15_io_to_pes_6_in_valid),
    .io_to_pes_6_in_bits(PENetwork_15_io_to_pes_6_in_bits),
    .io_to_pes_6_out_valid(PENetwork_15_io_to_pes_6_out_valid),
    .io_to_pes_6_out_bits(PENetwork_15_io_to_pes_6_out_bits),
    .io_to_pes_7_in_valid(PENetwork_15_io_to_pes_7_in_valid),
    .io_to_pes_7_in_bits(PENetwork_15_io_to_pes_7_in_bits),
    .io_to_pes_7_out_valid(PENetwork_15_io_to_pes_7_out_valid),
    .io_to_pes_7_out_bits(PENetwork_15_io_to_pes_7_out_bits),
    .io_to_mem_valid(PENetwork_15_io_to_mem_valid),
    .io_to_mem_bits(PENetwork_15_io_to_mem_bits)
  );
  PENetwork_16 PENetwork_16 ( // @[pearray.scala 134:13]
    .io_to_pes_0_in_valid(PENetwork_16_io_to_pes_0_in_valid),
    .io_to_pes_0_in_bits(PENetwork_16_io_to_pes_0_in_bits),
    .io_to_pes_0_out_valid(PENetwork_16_io_to_pes_0_out_valid),
    .io_to_pes_0_out_bits(PENetwork_16_io_to_pes_0_out_bits),
    .io_to_pes_1_in_valid(PENetwork_16_io_to_pes_1_in_valid),
    .io_to_pes_1_in_bits(PENetwork_16_io_to_pes_1_in_bits),
    .io_to_pes_1_out_valid(PENetwork_16_io_to_pes_1_out_valid),
    .io_to_pes_1_out_bits(PENetwork_16_io_to_pes_1_out_bits),
    .io_to_pes_2_in_valid(PENetwork_16_io_to_pes_2_in_valid),
    .io_to_pes_2_in_bits(PENetwork_16_io_to_pes_2_in_bits),
    .io_to_pes_2_out_valid(PENetwork_16_io_to_pes_2_out_valid),
    .io_to_pes_2_out_bits(PENetwork_16_io_to_pes_2_out_bits),
    .io_to_pes_3_in_valid(PENetwork_16_io_to_pes_3_in_valid),
    .io_to_pes_3_in_bits(PENetwork_16_io_to_pes_3_in_bits),
    .io_to_pes_3_out_valid(PENetwork_16_io_to_pes_3_out_valid),
    .io_to_pes_3_out_bits(PENetwork_16_io_to_pes_3_out_bits),
    .io_to_pes_4_in_valid(PENetwork_16_io_to_pes_4_in_valid),
    .io_to_pes_4_in_bits(PENetwork_16_io_to_pes_4_in_bits),
    .io_to_pes_4_out_valid(PENetwork_16_io_to_pes_4_out_valid),
    .io_to_pes_4_out_bits(PENetwork_16_io_to_pes_4_out_bits),
    .io_to_pes_5_in_valid(PENetwork_16_io_to_pes_5_in_valid),
    .io_to_pes_5_in_bits(PENetwork_16_io_to_pes_5_in_bits),
    .io_to_pes_5_out_valid(PENetwork_16_io_to_pes_5_out_valid),
    .io_to_pes_5_out_bits(PENetwork_16_io_to_pes_5_out_bits),
    .io_to_pes_6_in_valid(PENetwork_16_io_to_pes_6_in_valid),
    .io_to_pes_6_in_bits(PENetwork_16_io_to_pes_6_in_bits),
    .io_to_pes_6_out_valid(PENetwork_16_io_to_pes_6_out_valid),
    .io_to_pes_6_out_bits(PENetwork_16_io_to_pes_6_out_bits),
    .io_to_pes_7_in_valid(PENetwork_16_io_to_pes_7_in_valid),
    .io_to_pes_7_in_bits(PENetwork_16_io_to_pes_7_in_bits),
    .io_to_mem_valid(PENetwork_16_io_to_mem_valid),
    .io_to_mem_bits(PENetwork_16_io_to_mem_bits)
  );
  PENetwork_16 PENetwork_17 ( // @[pearray.scala 134:13]
    .io_to_pes_0_in_valid(PENetwork_17_io_to_pes_0_in_valid),
    .io_to_pes_0_in_bits(PENetwork_17_io_to_pes_0_in_bits),
    .io_to_pes_0_out_valid(PENetwork_17_io_to_pes_0_out_valid),
    .io_to_pes_0_out_bits(PENetwork_17_io_to_pes_0_out_bits),
    .io_to_pes_1_in_valid(PENetwork_17_io_to_pes_1_in_valid),
    .io_to_pes_1_in_bits(PENetwork_17_io_to_pes_1_in_bits),
    .io_to_pes_1_out_valid(PENetwork_17_io_to_pes_1_out_valid),
    .io_to_pes_1_out_bits(PENetwork_17_io_to_pes_1_out_bits),
    .io_to_pes_2_in_valid(PENetwork_17_io_to_pes_2_in_valid),
    .io_to_pes_2_in_bits(PENetwork_17_io_to_pes_2_in_bits),
    .io_to_pes_2_out_valid(PENetwork_17_io_to_pes_2_out_valid),
    .io_to_pes_2_out_bits(PENetwork_17_io_to_pes_2_out_bits),
    .io_to_pes_3_in_valid(PENetwork_17_io_to_pes_3_in_valid),
    .io_to_pes_3_in_bits(PENetwork_17_io_to_pes_3_in_bits),
    .io_to_pes_3_out_valid(PENetwork_17_io_to_pes_3_out_valid),
    .io_to_pes_3_out_bits(PENetwork_17_io_to_pes_3_out_bits),
    .io_to_pes_4_in_valid(PENetwork_17_io_to_pes_4_in_valid),
    .io_to_pes_4_in_bits(PENetwork_17_io_to_pes_4_in_bits),
    .io_to_pes_4_out_valid(PENetwork_17_io_to_pes_4_out_valid),
    .io_to_pes_4_out_bits(PENetwork_17_io_to_pes_4_out_bits),
    .io_to_pes_5_in_valid(PENetwork_17_io_to_pes_5_in_valid),
    .io_to_pes_5_in_bits(PENetwork_17_io_to_pes_5_in_bits),
    .io_to_pes_5_out_valid(PENetwork_17_io_to_pes_5_out_valid),
    .io_to_pes_5_out_bits(PENetwork_17_io_to_pes_5_out_bits),
    .io_to_pes_6_in_valid(PENetwork_17_io_to_pes_6_in_valid),
    .io_to_pes_6_in_bits(PENetwork_17_io_to_pes_6_in_bits),
    .io_to_pes_6_out_valid(PENetwork_17_io_to_pes_6_out_valid),
    .io_to_pes_6_out_bits(PENetwork_17_io_to_pes_6_out_bits),
    .io_to_pes_7_in_valid(PENetwork_17_io_to_pes_7_in_valid),
    .io_to_pes_7_in_bits(PENetwork_17_io_to_pes_7_in_bits),
    .io_to_mem_valid(PENetwork_17_io_to_mem_valid),
    .io_to_mem_bits(PENetwork_17_io_to_mem_bits)
  );
  PENetwork_16 PENetwork_18 ( // @[pearray.scala 134:13]
    .io_to_pes_0_in_valid(PENetwork_18_io_to_pes_0_in_valid),
    .io_to_pes_0_in_bits(PENetwork_18_io_to_pes_0_in_bits),
    .io_to_pes_0_out_valid(PENetwork_18_io_to_pes_0_out_valid),
    .io_to_pes_0_out_bits(PENetwork_18_io_to_pes_0_out_bits),
    .io_to_pes_1_in_valid(PENetwork_18_io_to_pes_1_in_valid),
    .io_to_pes_1_in_bits(PENetwork_18_io_to_pes_1_in_bits),
    .io_to_pes_1_out_valid(PENetwork_18_io_to_pes_1_out_valid),
    .io_to_pes_1_out_bits(PENetwork_18_io_to_pes_1_out_bits),
    .io_to_pes_2_in_valid(PENetwork_18_io_to_pes_2_in_valid),
    .io_to_pes_2_in_bits(PENetwork_18_io_to_pes_2_in_bits),
    .io_to_pes_2_out_valid(PENetwork_18_io_to_pes_2_out_valid),
    .io_to_pes_2_out_bits(PENetwork_18_io_to_pes_2_out_bits),
    .io_to_pes_3_in_valid(PENetwork_18_io_to_pes_3_in_valid),
    .io_to_pes_3_in_bits(PENetwork_18_io_to_pes_3_in_bits),
    .io_to_pes_3_out_valid(PENetwork_18_io_to_pes_3_out_valid),
    .io_to_pes_3_out_bits(PENetwork_18_io_to_pes_3_out_bits),
    .io_to_pes_4_in_valid(PENetwork_18_io_to_pes_4_in_valid),
    .io_to_pes_4_in_bits(PENetwork_18_io_to_pes_4_in_bits),
    .io_to_pes_4_out_valid(PENetwork_18_io_to_pes_4_out_valid),
    .io_to_pes_4_out_bits(PENetwork_18_io_to_pes_4_out_bits),
    .io_to_pes_5_in_valid(PENetwork_18_io_to_pes_5_in_valid),
    .io_to_pes_5_in_bits(PENetwork_18_io_to_pes_5_in_bits),
    .io_to_pes_5_out_valid(PENetwork_18_io_to_pes_5_out_valid),
    .io_to_pes_5_out_bits(PENetwork_18_io_to_pes_5_out_bits),
    .io_to_pes_6_in_valid(PENetwork_18_io_to_pes_6_in_valid),
    .io_to_pes_6_in_bits(PENetwork_18_io_to_pes_6_in_bits),
    .io_to_pes_6_out_valid(PENetwork_18_io_to_pes_6_out_valid),
    .io_to_pes_6_out_bits(PENetwork_18_io_to_pes_6_out_bits),
    .io_to_pes_7_in_valid(PENetwork_18_io_to_pes_7_in_valid),
    .io_to_pes_7_in_bits(PENetwork_18_io_to_pes_7_in_bits),
    .io_to_mem_valid(PENetwork_18_io_to_mem_valid),
    .io_to_mem_bits(PENetwork_18_io_to_mem_bits)
  );
  PENetwork_16 PENetwork_19 ( // @[pearray.scala 134:13]
    .io_to_pes_0_in_valid(PENetwork_19_io_to_pes_0_in_valid),
    .io_to_pes_0_in_bits(PENetwork_19_io_to_pes_0_in_bits),
    .io_to_pes_0_out_valid(PENetwork_19_io_to_pes_0_out_valid),
    .io_to_pes_0_out_bits(PENetwork_19_io_to_pes_0_out_bits),
    .io_to_pes_1_in_valid(PENetwork_19_io_to_pes_1_in_valid),
    .io_to_pes_1_in_bits(PENetwork_19_io_to_pes_1_in_bits),
    .io_to_pes_1_out_valid(PENetwork_19_io_to_pes_1_out_valid),
    .io_to_pes_1_out_bits(PENetwork_19_io_to_pes_1_out_bits),
    .io_to_pes_2_in_valid(PENetwork_19_io_to_pes_2_in_valid),
    .io_to_pes_2_in_bits(PENetwork_19_io_to_pes_2_in_bits),
    .io_to_pes_2_out_valid(PENetwork_19_io_to_pes_2_out_valid),
    .io_to_pes_2_out_bits(PENetwork_19_io_to_pes_2_out_bits),
    .io_to_pes_3_in_valid(PENetwork_19_io_to_pes_3_in_valid),
    .io_to_pes_3_in_bits(PENetwork_19_io_to_pes_3_in_bits),
    .io_to_pes_3_out_valid(PENetwork_19_io_to_pes_3_out_valid),
    .io_to_pes_3_out_bits(PENetwork_19_io_to_pes_3_out_bits),
    .io_to_pes_4_in_valid(PENetwork_19_io_to_pes_4_in_valid),
    .io_to_pes_4_in_bits(PENetwork_19_io_to_pes_4_in_bits),
    .io_to_pes_4_out_valid(PENetwork_19_io_to_pes_4_out_valid),
    .io_to_pes_4_out_bits(PENetwork_19_io_to_pes_4_out_bits),
    .io_to_pes_5_in_valid(PENetwork_19_io_to_pes_5_in_valid),
    .io_to_pes_5_in_bits(PENetwork_19_io_to_pes_5_in_bits),
    .io_to_pes_5_out_valid(PENetwork_19_io_to_pes_5_out_valid),
    .io_to_pes_5_out_bits(PENetwork_19_io_to_pes_5_out_bits),
    .io_to_pes_6_in_valid(PENetwork_19_io_to_pes_6_in_valid),
    .io_to_pes_6_in_bits(PENetwork_19_io_to_pes_6_in_bits),
    .io_to_pes_6_out_valid(PENetwork_19_io_to_pes_6_out_valid),
    .io_to_pes_6_out_bits(PENetwork_19_io_to_pes_6_out_bits),
    .io_to_pes_7_in_valid(PENetwork_19_io_to_pes_7_in_valid),
    .io_to_pes_7_in_bits(PENetwork_19_io_to_pes_7_in_bits),
    .io_to_mem_valid(PENetwork_19_io_to_mem_valid),
    .io_to_mem_bits(PENetwork_19_io_to_mem_bits)
  );
  PENetwork_16 PENetwork_20 ( // @[pearray.scala 134:13]
    .io_to_pes_0_in_valid(PENetwork_20_io_to_pes_0_in_valid),
    .io_to_pes_0_in_bits(PENetwork_20_io_to_pes_0_in_bits),
    .io_to_pes_0_out_valid(PENetwork_20_io_to_pes_0_out_valid),
    .io_to_pes_0_out_bits(PENetwork_20_io_to_pes_0_out_bits),
    .io_to_pes_1_in_valid(PENetwork_20_io_to_pes_1_in_valid),
    .io_to_pes_1_in_bits(PENetwork_20_io_to_pes_1_in_bits),
    .io_to_pes_1_out_valid(PENetwork_20_io_to_pes_1_out_valid),
    .io_to_pes_1_out_bits(PENetwork_20_io_to_pes_1_out_bits),
    .io_to_pes_2_in_valid(PENetwork_20_io_to_pes_2_in_valid),
    .io_to_pes_2_in_bits(PENetwork_20_io_to_pes_2_in_bits),
    .io_to_pes_2_out_valid(PENetwork_20_io_to_pes_2_out_valid),
    .io_to_pes_2_out_bits(PENetwork_20_io_to_pes_2_out_bits),
    .io_to_pes_3_in_valid(PENetwork_20_io_to_pes_3_in_valid),
    .io_to_pes_3_in_bits(PENetwork_20_io_to_pes_3_in_bits),
    .io_to_pes_3_out_valid(PENetwork_20_io_to_pes_3_out_valid),
    .io_to_pes_3_out_bits(PENetwork_20_io_to_pes_3_out_bits),
    .io_to_pes_4_in_valid(PENetwork_20_io_to_pes_4_in_valid),
    .io_to_pes_4_in_bits(PENetwork_20_io_to_pes_4_in_bits),
    .io_to_pes_4_out_valid(PENetwork_20_io_to_pes_4_out_valid),
    .io_to_pes_4_out_bits(PENetwork_20_io_to_pes_4_out_bits),
    .io_to_pes_5_in_valid(PENetwork_20_io_to_pes_5_in_valid),
    .io_to_pes_5_in_bits(PENetwork_20_io_to_pes_5_in_bits),
    .io_to_pes_5_out_valid(PENetwork_20_io_to_pes_5_out_valid),
    .io_to_pes_5_out_bits(PENetwork_20_io_to_pes_5_out_bits),
    .io_to_pes_6_in_valid(PENetwork_20_io_to_pes_6_in_valid),
    .io_to_pes_6_in_bits(PENetwork_20_io_to_pes_6_in_bits),
    .io_to_pes_6_out_valid(PENetwork_20_io_to_pes_6_out_valid),
    .io_to_pes_6_out_bits(PENetwork_20_io_to_pes_6_out_bits),
    .io_to_pes_7_in_valid(PENetwork_20_io_to_pes_7_in_valid),
    .io_to_pes_7_in_bits(PENetwork_20_io_to_pes_7_in_bits),
    .io_to_mem_valid(PENetwork_20_io_to_mem_valid),
    .io_to_mem_bits(PENetwork_20_io_to_mem_bits)
  );
  PENetwork_16 PENetwork_21 ( // @[pearray.scala 134:13]
    .io_to_pes_0_in_valid(PENetwork_21_io_to_pes_0_in_valid),
    .io_to_pes_0_in_bits(PENetwork_21_io_to_pes_0_in_bits),
    .io_to_pes_0_out_valid(PENetwork_21_io_to_pes_0_out_valid),
    .io_to_pes_0_out_bits(PENetwork_21_io_to_pes_0_out_bits),
    .io_to_pes_1_in_valid(PENetwork_21_io_to_pes_1_in_valid),
    .io_to_pes_1_in_bits(PENetwork_21_io_to_pes_1_in_bits),
    .io_to_pes_1_out_valid(PENetwork_21_io_to_pes_1_out_valid),
    .io_to_pes_1_out_bits(PENetwork_21_io_to_pes_1_out_bits),
    .io_to_pes_2_in_valid(PENetwork_21_io_to_pes_2_in_valid),
    .io_to_pes_2_in_bits(PENetwork_21_io_to_pes_2_in_bits),
    .io_to_pes_2_out_valid(PENetwork_21_io_to_pes_2_out_valid),
    .io_to_pes_2_out_bits(PENetwork_21_io_to_pes_2_out_bits),
    .io_to_pes_3_in_valid(PENetwork_21_io_to_pes_3_in_valid),
    .io_to_pes_3_in_bits(PENetwork_21_io_to_pes_3_in_bits),
    .io_to_pes_3_out_valid(PENetwork_21_io_to_pes_3_out_valid),
    .io_to_pes_3_out_bits(PENetwork_21_io_to_pes_3_out_bits),
    .io_to_pes_4_in_valid(PENetwork_21_io_to_pes_4_in_valid),
    .io_to_pes_4_in_bits(PENetwork_21_io_to_pes_4_in_bits),
    .io_to_pes_4_out_valid(PENetwork_21_io_to_pes_4_out_valid),
    .io_to_pes_4_out_bits(PENetwork_21_io_to_pes_4_out_bits),
    .io_to_pes_5_in_valid(PENetwork_21_io_to_pes_5_in_valid),
    .io_to_pes_5_in_bits(PENetwork_21_io_to_pes_5_in_bits),
    .io_to_pes_5_out_valid(PENetwork_21_io_to_pes_5_out_valid),
    .io_to_pes_5_out_bits(PENetwork_21_io_to_pes_5_out_bits),
    .io_to_pes_6_in_valid(PENetwork_21_io_to_pes_6_in_valid),
    .io_to_pes_6_in_bits(PENetwork_21_io_to_pes_6_in_bits),
    .io_to_pes_6_out_valid(PENetwork_21_io_to_pes_6_out_valid),
    .io_to_pes_6_out_bits(PENetwork_21_io_to_pes_6_out_bits),
    .io_to_pes_7_in_valid(PENetwork_21_io_to_pes_7_in_valid),
    .io_to_pes_7_in_bits(PENetwork_21_io_to_pes_7_in_bits),
    .io_to_mem_valid(PENetwork_21_io_to_mem_valid),
    .io_to_mem_bits(PENetwork_21_io_to_mem_bits)
  );
  PENetwork_16 PENetwork_22 ( // @[pearray.scala 134:13]
    .io_to_pes_0_in_valid(PENetwork_22_io_to_pes_0_in_valid),
    .io_to_pes_0_in_bits(PENetwork_22_io_to_pes_0_in_bits),
    .io_to_pes_0_out_valid(PENetwork_22_io_to_pes_0_out_valid),
    .io_to_pes_0_out_bits(PENetwork_22_io_to_pes_0_out_bits),
    .io_to_pes_1_in_valid(PENetwork_22_io_to_pes_1_in_valid),
    .io_to_pes_1_in_bits(PENetwork_22_io_to_pes_1_in_bits),
    .io_to_pes_1_out_valid(PENetwork_22_io_to_pes_1_out_valid),
    .io_to_pes_1_out_bits(PENetwork_22_io_to_pes_1_out_bits),
    .io_to_pes_2_in_valid(PENetwork_22_io_to_pes_2_in_valid),
    .io_to_pes_2_in_bits(PENetwork_22_io_to_pes_2_in_bits),
    .io_to_pes_2_out_valid(PENetwork_22_io_to_pes_2_out_valid),
    .io_to_pes_2_out_bits(PENetwork_22_io_to_pes_2_out_bits),
    .io_to_pes_3_in_valid(PENetwork_22_io_to_pes_3_in_valid),
    .io_to_pes_3_in_bits(PENetwork_22_io_to_pes_3_in_bits),
    .io_to_pes_3_out_valid(PENetwork_22_io_to_pes_3_out_valid),
    .io_to_pes_3_out_bits(PENetwork_22_io_to_pes_3_out_bits),
    .io_to_pes_4_in_valid(PENetwork_22_io_to_pes_4_in_valid),
    .io_to_pes_4_in_bits(PENetwork_22_io_to_pes_4_in_bits),
    .io_to_pes_4_out_valid(PENetwork_22_io_to_pes_4_out_valid),
    .io_to_pes_4_out_bits(PENetwork_22_io_to_pes_4_out_bits),
    .io_to_pes_5_in_valid(PENetwork_22_io_to_pes_5_in_valid),
    .io_to_pes_5_in_bits(PENetwork_22_io_to_pes_5_in_bits),
    .io_to_pes_5_out_valid(PENetwork_22_io_to_pes_5_out_valid),
    .io_to_pes_5_out_bits(PENetwork_22_io_to_pes_5_out_bits),
    .io_to_pes_6_in_valid(PENetwork_22_io_to_pes_6_in_valid),
    .io_to_pes_6_in_bits(PENetwork_22_io_to_pes_6_in_bits),
    .io_to_pes_6_out_valid(PENetwork_22_io_to_pes_6_out_valid),
    .io_to_pes_6_out_bits(PENetwork_22_io_to_pes_6_out_bits),
    .io_to_pes_7_in_valid(PENetwork_22_io_to_pes_7_in_valid),
    .io_to_pes_7_in_bits(PENetwork_22_io_to_pes_7_in_bits),
    .io_to_mem_valid(PENetwork_22_io_to_mem_valid),
    .io_to_mem_bits(PENetwork_22_io_to_mem_bits)
  );
  PENetwork_16 PENetwork_23 ( // @[pearray.scala 134:13]
    .io_to_pes_0_in_valid(PENetwork_23_io_to_pes_0_in_valid),
    .io_to_pes_0_in_bits(PENetwork_23_io_to_pes_0_in_bits),
    .io_to_pes_0_out_valid(PENetwork_23_io_to_pes_0_out_valid),
    .io_to_pes_0_out_bits(PENetwork_23_io_to_pes_0_out_bits),
    .io_to_pes_1_in_valid(PENetwork_23_io_to_pes_1_in_valid),
    .io_to_pes_1_in_bits(PENetwork_23_io_to_pes_1_in_bits),
    .io_to_pes_1_out_valid(PENetwork_23_io_to_pes_1_out_valid),
    .io_to_pes_1_out_bits(PENetwork_23_io_to_pes_1_out_bits),
    .io_to_pes_2_in_valid(PENetwork_23_io_to_pes_2_in_valid),
    .io_to_pes_2_in_bits(PENetwork_23_io_to_pes_2_in_bits),
    .io_to_pes_2_out_valid(PENetwork_23_io_to_pes_2_out_valid),
    .io_to_pes_2_out_bits(PENetwork_23_io_to_pes_2_out_bits),
    .io_to_pes_3_in_valid(PENetwork_23_io_to_pes_3_in_valid),
    .io_to_pes_3_in_bits(PENetwork_23_io_to_pes_3_in_bits),
    .io_to_pes_3_out_valid(PENetwork_23_io_to_pes_3_out_valid),
    .io_to_pes_3_out_bits(PENetwork_23_io_to_pes_3_out_bits),
    .io_to_pes_4_in_valid(PENetwork_23_io_to_pes_4_in_valid),
    .io_to_pes_4_in_bits(PENetwork_23_io_to_pes_4_in_bits),
    .io_to_pes_4_out_valid(PENetwork_23_io_to_pes_4_out_valid),
    .io_to_pes_4_out_bits(PENetwork_23_io_to_pes_4_out_bits),
    .io_to_pes_5_in_valid(PENetwork_23_io_to_pes_5_in_valid),
    .io_to_pes_5_in_bits(PENetwork_23_io_to_pes_5_in_bits),
    .io_to_pes_5_out_valid(PENetwork_23_io_to_pes_5_out_valid),
    .io_to_pes_5_out_bits(PENetwork_23_io_to_pes_5_out_bits),
    .io_to_pes_6_in_valid(PENetwork_23_io_to_pes_6_in_valid),
    .io_to_pes_6_in_bits(PENetwork_23_io_to_pes_6_in_bits),
    .io_to_pes_6_out_valid(PENetwork_23_io_to_pes_6_out_valid),
    .io_to_pes_6_out_bits(PENetwork_23_io_to_pes_6_out_bits),
    .io_to_pes_7_in_valid(PENetwork_23_io_to_pes_7_in_valid),
    .io_to_pes_7_in_bits(PENetwork_23_io_to_pes_7_in_bits),
    .io_to_mem_valid(PENetwork_23_io_to_mem_valid),
    .io_to_mem_bits(PENetwork_23_io_to_mem_bits)
  );
  PENetwork_16 PENetwork_24 ( // @[pearray.scala 134:13]
    .io_to_pes_0_in_valid(PENetwork_24_io_to_pes_0_in_valid),
    .io_to_pes_0_in_bits(PENetwork_24_io_to_pes_0_in_bits),
    .io_to_pes_0_out_valid(PENetwork_24_io_to_pes_0_out_valid),
    .io_to_pes_0_out_bits(PENetwork_24_io_to_pes_0_out_bits),
    .io_to_pes_1_in_valid(PENetwork_24_io_to_pes_1_in_valid),
    .io_to_pes_1_in_bits(PENetwork_24_io_to_pes_1_in_bits),
    .io_to_pes_1_out_valid(PENetwork_24_io_to_pes_1_out_valid),
    .io_to_pes_1_out_bits(PENetwork_24_io_to_pes_1_out_bits),
    .io_to_pes_2_in_valid(PENetwork_24_io_to_pes_2_in_valid),
    .io_to_pes_2_in_bits(PENetwork_24_io_to_pes_2_in_bits),
    .io_to_pes_2_out_valid(PENetwork_24_io_to_pes_2_out_valid),
    .io_to_pes_2_out_bits(PENetwork_24_io_to_pes_2_out_bits),
    .io_to_pes_3_in_valid(PENetwork_24_io_to_pes_3_in_valid),
    .io_to_pes_3_in_bits(PENetwork_24_io_to_pes_3_in_bits),
    .io_to_pes_3_out_valid(PENetwork_24_io_to_pes_3_out_valid),
    .io_to_pes_3_out_bits(PENetwork_24_io_to_pes_3_out_bits),
    .io_to_pes_4_in_valid(PENetwork_24_io_to_pes_4_in_valid),
    .io_to_pes_4_in_bits(PENetwork_24_io_to_pes_4_in_bits),
    .io_to_pes_4_out_valid(PENetwork_24_io_to_pes_4_out_valid),
    .io_to_pes_4_out_bits(PENetwork_24_io_to_pes_4_out_bits),
    .io_to_pes_5_in_valid(PENetwork_24_io_to_pes_5_in_valid),
    .io_to_pes_5_in_bits(PENetwork_24_io_to_pes_5_in_bits),
    .io_to_pes_5_out_valid(PENetwork_24_io_to_pes_5_out_valid),
    .io_to_pes_5_out_bits(PENetwork_24_io_to_pes_5_out_bits),
    .io_to_pes_6_in_valid(PENetwork_24_io_to_pes_6_in_valid),
    .io_to_pes_6_in_bits(PENetwork_24_io_to_pes_6_in_bits),
    .io_to_pes_6_out_valid(PENetwork_24_io_to_pes_6_out_valid),
    .io_to_pes_6_out_bits(PENetwork_24_io_to_pes_6_out_bits),
    .io_to_pes_7_in_valid(PENetwork_24_io_to_pes_7_in_valid),
    .io_to_pes_7_in_bits(PENetwork_24_io_to_pes_7_in_bits),
    .io_to_mem_valid(PENetwork_24_io_to_mem_valid),
    .io_to_mem_bits(PENetwork_24_io_to_mem_bits)
  );
  PENetwork_16 PENetwork_25 ( // @[pearray.scala 134:13]
    .io_to_pes_0_in_valid(PENetwork_25_io_to_pes_0_in_valid),
    .io_to_pes_0_in_bits(PENetwork_25_io_to_pes_0_in_bits),
    .io_to_pes_0_out_valid(PENetwork_25_io_to_pes_0_out_valid),
    .io_to_pes_0_out_bits(PENetwork_25_io_to_pes_0_out_bits),
    .io_to_pes_1_in_valid(PENetwork_25_io_to_pes_1_in_valid),
    .io_to_pes_1_in_bits(PENetwork_25_io_to_pes_1_in_bits),
    .io_to_pes_1_out_valid(PENetwork_25_io_to_pes_1_out_valid),
    .io_to_pes_1_out_bits(PENetwork_25_io_to_pes_1_out_bits),
    .io_to_pes_2_in_valid(PENetwork_25_io_to_pes_2_in_valid),
    .io_to_pes_2_in_bits(PENetwork_25_io_to_pes_2_in_bits),
    .io_to_pes_2_out_valid(PENetwork_25_io_to_pes_2_out_valid),
    .io_to_pes_2_out_bits(PENetwork_25_io_to_pes_2_out_bits),
    .io_to_pes_3_in_valid(PENetwork_25_io_to_pes_3_in_valid),
    .io_to_pes_3_in_bits(PENetwork_25_io_to_pes_3_in_bits),
    .io_to_pes_3_out_valid(PENetwork_25_io_to_pes_3_out_valid),
    .io_to_pes_3_out_bits(PENetwork_25_io_to_pes_3_out_bits),
    .io_to_pes_4_in_valid(PENetwork_25_io_to_pes_4_in_valid),
    .io_to_pes_4_in_bits(PENetwork_25_io_to_pes_4_in_bits),
    .io_to_pes_4_out_valid(PENetwork_25_io_to_pes_4_out_valid),
    .io_to_pes_4_out_bits(PENetwork_25_io_to_pes_4_out_bits),
    .io_to_pes_5_in_valid(PENetwork_25_io_to_pes_5_in_valid),
    .io_to_pes_5_in_bits(PENetwork_25_io_to_pes_5_in_bits),
    .io_to_pes_5_out_valid(PENetwork_25_io_to_pes_5_out_valid),
    .io_to_pes_5_out_bits(PENetwork_25_io_to_pes_5_out_bits),
    .io_to_pes_6_in_valid(PENetwork_25_io_to_pes_6_in_valid),
    .io_to_pes_6_in_bits(PENetwork_25_io_to_pes_6_in_bits),
    .io_to_pes_6_out_valid(PENetwork_25_io_to_pes_6_out_valid),
    .io_to_pes_6_out_bits(PENetwork_25_io_to_pes_6_out_bits),
    .io_to_pes_7_in_valid(PENetwork_25_io_to_pes_7_in_valid),
    .io_to_pes_7_in_bits(PENetwork_25_io_to_pes_7_in_bits),
    .io_to_mem_valid(PENetwork_25_io_to_mem_valid),
    .io_to_mem_bits(PENetwork_25_io_to_mem_bits)
  );
  PENetwork_16 PENetwork_26 ( // @[pearray.scala 134:13]
    .io_to_pes_0_in_valid(PENetwork_26_io_to_pes_0_in_valid),
    .io_to_pes_0_in_bits(PENetwork_26_io_to_pes_0_in_bits),
    .io_to_pes_0_out_valid(PENetwork_26_io_to_pes_0_out_valid),
    .io_to_pes_0_out_bits(PENetwork_26_io_to_pes_0_out_bits),
    .io_to_pes_1_in_valid(PENetwork_26_io_to_pes_1_in_valid),
    .io_to_pes_1_in_bits(PENetwork_26_io_to_pes_1_in_bits),
    .io_to_pes_1_out_valid(PENetwork_26_io_to_pes_1_out_valid),
    .io_to_pes_1_out_bits(PENetwork_26_io_to_pes_1_out_bits),
    .io_to_pes_2_in_valid(PENetwork_26_io_to_pes_2_in_valid),
    .io_to_pes_2_in_bits(PENetwork_26_io_to_pes_2_in_bits),
    .io_to_pes_2_out_valid(PENetwork_26_io_to_pes_2_out_valid),
    .io_to_pes_2_out_bits(PENetwork_26_io_to_pes_2_out_bits),
    .io_to_pes_3_in_valid(PENetwork_26_io_to_pes_3_in_valid),
    .io_to_pes_3_in_bits(PENetwork_26_io_to_pes_3_in_bits),
    .io_to_pes_3_out_valid(PENetwork_26_io_to_pes_3_out_valid),
    .io_to_pes_3_out_bits(PENetwork_26_io_to_pes_3_out_bits),
    .io_to_pes_4_in_valid(PENetwork_26_io_to_pes_4_in_valid),
    .io_to_pes_4_in_bits(PENetwork_26_io_to_pes_4_in_bits),
    .io_to_pes_4_out_valid(PENetwork_26_io_to_pes_4_out_valid),
    .io_to_pes_4_out_bits(PENetwork_26_io_to_pes_4_out_bits),
    .io_to_pes_5_in_valid(PENetwork_26_io_to_pes_5_in_valid),
    .io_to_pes_5_in_bits(PENetwork_26_io_to_pes_5_in_bits),
    .io_to_pes_5_out_valid(PENetwork_26_io_to_pes_5_out_valid),
    .io_to_pes_5_out_bits(PENetwork_26_io_to_pes_5_out_bits),
    .io_to_pes_6_in_valid(PENetwork_26_io_to_pes_6_in_valid),
    .io_to_pes_6_in_bits(PENetwork_26_io_to_pes_6_in_bits),
    .io_to_pes_6_out_valid(PENetwork_26_io_to_pes_6_out_valid),
    .io_to_pes_6_out_bits(PENetwork_26_io_to_pes_6_out_bits),
    .io_to_pes_7_in_valid(PENetwork_26_io_to_pes_7_in_valid),
    .io_to_pes_7_in_bits(PENetwork_26_io_to_pes_7_in_bits),
    .io_to_mem_valid(PENetwork_26_io_to_mem_valid),
    .io_to_mem_bits(PENetwork_26_io_to_mem_bits)
  );
  PENetwork_16 PENetwork_27 ( // @[pearray.scala 134:13]
    .io_to_pes_0_in_valid(PENetwork_27_io_to_pes_0_in_valid),
    .io_to_pes_0_in_bits(PENetwork_27_io_to_pes_0_in_bits),
    .io_to_pes_0_out_valid(PENetwork_27_io_to_pes_0_out_valid),
    .io_to_pes_0_out_bits(PENetwork_27_io_to_pes_0_out_bits),
    .io_to_pes_1_in_valid(PENetwork_27_io_to_pes_1_in_valid),
    .io_to_pes_1_in_bits(PENetwork_27_io_to_pes_1_in_bits),
    .io_to_pes_1_out_valid(PENetwork_27_io_to_pes_1_out_valid),
    .io_to_pes_1_out_bits(PENetwork_27_io_to_pes_1_out_bits),
    .io_to_pes_2_in_valid(PENetwork_27_io_to_pes_2_in_valid),
    .io_to_pes_2_in_bits(PENetwork_27_io_to_pes_2_in_bits),
    .io_to_pes_2_out_valid(PENetwork_27_io_to_pes_2_out_valid),
    .io_to_pes_2_out_bits(PENetwork_27_io_to_pes_2_out_bits),
    .io_to_pes_3_in_valid(PENetwork_27_io_to_pes_3_in_valid),
    .io_to_pes_3_in_bits(PENetwork_27_io_to_pes_3_in_bits),
    .io_to_pes_3_out_valid(PENetwork_27_io_to_pes_3_out_valid),
    .io_to_pes_3_out_bits(PENetwork_27_io_to_pes_3_out_bits),
    .io_to_pes_4_in_valid(PENetwork_27_io_to_pes_4_in_valid),
    .io_to_pes_4_in_bits(PENetwork_27_io_to_pes_4_in_bits),
    .io_to_pes_4_out_valid(PENetwork_27_io_to_pes_4_out_valid),
    .io_to_pes_4_out_bits(PENetwork_27_io_to_pes_4_out_bits),
    .io_to_pes_5_in_valid(PENetwork_27_io_to_pes_5_in_valid),
    .io_to_pes_5_in_bits(PENetwork_27_io_to_pes_5_in_bits),
    .io_to_pes_5_out_valid(PENetwork_27_io_to_pes_5_out_valid),
    .io_to_pes_5_out_bits(PENetwork_27_io_to_pes_5_out_bits),
    .io_to_pes_6_in_valid(PENetwork_27_io_to_pes_6_in_valid),
    .io_to_pes_6_in_bits(PENetwork_27_io_to_pes_6_in_bits),
    .io_to_pes_6_out_valid(PENetwork_27_io_to_pes_6_out_valid),
    .io_to_pes_6_out_bits(PENetwork_27_io_to_pes_6_out_bits),
    .io_to_pes_7_in_valid(PENetwork_27_io_to_pes_7_in_valid),
    .io_to_pes_7_in_bits(PENetwork_27_io_to_pes_7_in_bits),
    .io_to_mem_valid(PENetwork_27_io_to_mem_valid),
    .io_to_mem_bits(PENetwork_27_io_to_mem_bits)
  );
  PENetwork_16 PENetwork_28 ( // @[pearray.scala 134:13]
    .io_to_pes_0_in_valid(PENetwork_28_io_to_pes_0_in_valid),
    .io_to_pes_0_in_bits(PENetwork_28_io_to_pes_0_in_bits),
    .io_to_pes_0_out_valid(PENetwork_28_io_to_pes_0_out_valid),
    .io_to_pes_0_out_bits(PENetwork_28_io_to_pes_0_out_bits),
    .io_to_pes_1_in_valid(PENetwork_28_io_to_pes_1_in_valid),
    .io_to_pes_1_in_bits(PENetwork_28_io_to_pes_1_in_bits),
    .io_to_pes_1_out_valid(PENetwork_28_io_to_pes_1_out_valid),
    .io_to_pes_1_out_bits(PENetwork_28_io_to_pes_1_out_bits),
    .io_to_pes_2_in_valid(PENetwork_28_io_to_pes_2_in_valid),
    .io_to_pes_2_in_bits(PENetwork_28_io_to_pes_2_in_bits),
    .io_to_pes_2_out_valid(PENetwork_28_io_to_pes_2_out_valid),
    .io_to_pes_2_out_bits(PENetwork_28_io_to_pes_2_out_bits),
    .io_to_pes_3_in_valid(PENetwork_28_io_to_pes_3_in_valid),
    .io_to_pes_3_in_bits(PENetwork_28_io_to_pes_3_in_bits),
    .io_to_pes_3_out_valid(PENetwork_28_io_to_pes_3_out_valid),
    .io_to_pes_3_out_bits(PENetwork_28_io_to_pes_3_out_bits),
    .io_to_pes_4_in_valid(PENetwork_28_io_to_pes_4_in_valid),
    .io_to_pes_4_in_bits(PENetwork_28_io_to_pes_4_in_bits),
    .io_to_pes_4_out_valid(PENetwork_28_io_to_pes_4_out_valid),
    .io_to_pes_4_out_bits(PENetwork_28_io_to_pes_4_out_bits),
    .io_to_pes_5_in_valid(PENetwork_28_io_to_pes_5_in_valid),
    .io_to_pes_5_in_bits(PENetwork_28_io_to_pes_5_in_bits),
    .io_to_pes_5_out_valid(PENetwork_28_io_to_pes_5_out_valid),
    .io_to_pes_5_out_bits(PENetwork_28_io_to_pes_5_out_bits),
    .io_to_pes_6_in_valid(PENetwork_28_io_to_pes_6_in_valid),
    .io_to_pes_6_in_bits(PENetwork_28_io_to_pes_6_in_bits),
    .io_to_pes_6_out_valid(PENetwork_28_io_to_pes_6_out_valid),
    .io_to_pes_6_out_bits(PENetwork_28_io_to_pes_6_out_bits),
    .io_to_pes_7_in_valid(PENetwork_28_io_to_pes_7_in_valid),
    .io_to_pes_7_in_bits(PENetwork_28_io_to_pes_7_in_bits),
    .io_to_mem_valid(PENetwork_28_io_to_mem_valid),
    .io_to_mem_bits(PENetwork_28_io_to_mem_bits)
  );
  PENetwork_16 PENetwork_29 ( // @[pearray.scala 134:13]
    .io_to_pes_0_in_valid(PENetwork_29_io_to_pes_0_in_valid),
    .io_to_pes_0_in_bits(PENetwork_29_io_to_pes_0_in_bits),
    .io_to_pes_0_out_valid(PENetwork_29_io_to_pes_0_out_valid),
    .io_to_pes_0_out_bits(PENetwork_29_io_to_pes_0_out_bits),
    .io_to_pes_1_in_valid(PENetwork_29_io_to_pes_1_in_valid),
    .io_to_pes_1_in_bits(PENetwork_29_io_to_pes_1_in_bits),
    .io_to_pes_1_out_valid(PENetwork_29_io_to_pes_1_out_valid),
    .io_to_pes_1_out_bits(PENetwork_29_io_to_pes_1_out_bits),
    .io_to_pes_2_in_valid(PENetwork_29_io_to_pes_2_in_valid),
    .io_to_pes_2_in_bits(PENetwork_29_io_to_pes_2_in_bits),
    .io_to_pes_2_out_valid(PENetwork_29_io_to_pes_2_out_valid),
    .io_to_pes_2_out_bits(PENetwork_29_io_to_pes_2_out_bits),
    .io_to_pes_3_in_valid(PENetwork_29_io_to_pes_3_in_valid),
    .io_to_pes_3_in_bits(PENetwork_29_io_to_pes_3_in_bits),
    .io_to_pes_3_out_valid(PENetwork_29_io_to_pes_3_out_valid),
    .io_to_pes_3_out_bits(PENetwork_29_io_to_pes_3_out_bits),
    .io_to_pes_4_in_valid(PENetwork_29_io_to_pes_4_in_valid),
    .io_to_pes_4_in_bits(PENetwork_29_io_to_pes_4_in_bits),
    .io_to_pes_4_out_valid(PENetwork_29_io_to_pes_4_out_valid),
    .io_to_pes_4_out_bits(PENetwork_29_io_to_pes_4_out_bits),
    .io_to_pes_5_in_valid(PENetwork_29_io_to_pes_5_in_valid),
    .io_to_pes_5_in_bits(PENetwork_29_io_to_pes_5_in_bits),
    .io_to_pes_5_out_valid(PENetwork_29_io_to_pes_5_out_valid),
    .io_to_pes_5_out_bits(PENetwork_29_io_to_pes_5_out_bits),
    .io_to_pes_6_in_valid(PENetwork_29_io_to_pes_6_in_valid),
    .io_to_pes_6_in_bits(PENetwork_29_io_to_pes_6_in_bits),
    .io_to_pes_6_out_valid(PENetwork_29_io_to_pes_6_out_valid),
    .io_to_pes_6_out_bits(PENetwork_29_io_to_pes_6_out_bits),
    .io_to_pes_7_in_valid(PENetwork_29_io_to_pes_7_in_valid),
    .io_to_pes_7_in_bits(PENetwork_29_io_to_pes_7_in_bits),
    .io_to_mem_valid(PENetwork_29_io_to_mem_valid),
    .io_to_mem_bits(PENetwork_29_io_to_mem_bits)
  );
  PENetwork_16 PENetwork_30 ( // @[pearray.scala 134:13]
    .io_to_pes_0_in_valid(PENetwork_30_io_to_pes_0_in_valid),
    .io_to_pes_0_in_bits(PENetwork_30_io_to_pes_0_in_bits),
    .io_to_pes_0_out_valid(PENetwork_30_io_to_pes_0_out_valid),
    .io_to_pes_0_out_bits(PENetwork_30_io_to_pes_0_out_bits),
    .io_to_pes_1_in_valid(PENetwork_30_io_to_pes_1_in_valid),
    .io_to_pes_1_in_bits(PENetwork_30_io_to_pes_1_in_bits),
    .io_to_pes_1_out_valid(PENetwork_30_io_to_pes_1_out_valid),
    .io_to_pes_1_out_bits(PENetwork_30_io_to_pes_1_out_bits),
    .io_to_pes_2_in_valid(PENetwork_30_io_to_pes_2_in_valid),
    .io_to_pes_2_in_bits(PENetwork_30_io_to_pes_2_in_bits),
    .io_to_pes_2_out_valid(PENetwork_30_io_to_pes_2_out_valid),
    .io_to_pes_2_out_bits(PENetwork_30_io_to_pes_2_out_bits),
    .io_to_pes_3_in_valid(PENetwork_30_io_to_pes_3_in_valid),
    .io_to_pes_3_in_bits(PENetwork_30_io_to_pes_3_in_bits),
    .io_to_pes_3_out_valid(PENetwork_30_io_to_pes_3_out_valid),
    .io_to_pes_3_out_bits(PENetwork_30_io_to_pes_3_out_bits),
    .io_to_pes_4_in_valid(PENetwork_30_io_to_pes_4_in_valid),
    .io_to_pes_4_in_bits(PENetwork_30_io_to_pes_4_in_bits),
    .io_to_pes_4_out_valid(PENetwork_30_io_to_pes_4_out_valid),
    .io_to_pes_4_out_bits(PENetwork_30_io_to_pes_4_out_bits),
    .io_to_pes_5_in_valid(PENetwork_30_io_to_pes_5_in_valid),
    .io_to_pes_5_in_bits(PENetwork_30_io_to_pes_5_in_bits),
    .io_to_pes_5_out_valid(PENetwork_30_io_to_pes_5_out_valid),
    .io_to_pes_5_out_bits(PENetwork_30_io_to_pes_5_out_bits),
    .io_to_pes_6_in_valid(PENetwork_30_io_to_pes_6_in_valid),
    .io_to_pes_6_in_bits(PENetwork_30_io_to_pes_6_in_bits),
    .io_to_pes_6_out_valid(PENetwork_30_io_to_pes_6_out_valid),
    .io_to_pes_6_out_bits(PENetwork_30_io_to_pes_6_out_bits),
    .io_to_pes_7_in_valid(PENetwork_30_io_to_pes_7_in_valid),
    .io_to_pes_7_in_bits(PENetwork_30_io_to_pes_7_in_bits),
    .io_to_mem_valid(PENetwork_30_io_to_mem_valid),
    .io_to_mem_bits(PENetwork_30_io_to_mem_bits)
  );
  PENetwork_16 PENetwork_31 ( // @[pearray.scala 134:13]
    .io_to_pes_0_in_valid(PENetwork_31_io_to_pes_0_in_valid),
    .io_to_pes_0_in_bits(PENetwork_31_io_to_pes_0_in_bits),
    .io_to_pes_0_out_valid(PENetwork_31_io_to_pes_0_out_valid),
    .io_to_pes_0_out_bits(PENetwork_31_io_to_pes_0_out_bits),
    .io_to_pes_1_in_valid(PENetwork_31_io_to_pes_1_in_valid),
    .io_to_pes_1_in_bits(PENetwork_31_io_to_pes_1_in_bits),
    .io_to_pes_1_out_valid(PENetwork_31_io_to_pes_1_out_valid),
    .io_to_pes_1_out_bits(PENetwork_31_io_to_pes_1_out_bits),
    .io_to_pes_2_in_valid(PENetwork_31_io_to_pes_2_in_valid),
    .io_to_pes_2_in_bits(PENetwork_31_io_to_pes_2_in_bits),
    .io_to_pes_2_out_valid(PENetwork_31_io_to_pes_2_out_valid),
    .io_to_pes_2_out_bits(PENetwork_31_io_to_pes_2_out_bits),
    .io_to_pes_3_in_valid(PENetwork_31_io_to_pes_3_in_valid),
    .io_to_pes_3_in_bits(PENetwork_31_io_to_pes_3_in_bits),
    .io_to_pes_3_out_valid(PENetwork_31_io_to_pes_3_out_valid),
    .io_to_pes_3_out_bits(PENetwork_31_io_to_pes_3_out_bits),
    .io_to_pes_4_in_valid(PENetwork_31_io_to_pes_4_in_valid),
    .io_to_pes_4_in_bits(PENetwork_31_io_to_pes_4_in_bits),
    .io_to_pes_4_out_valid(PENetwork_31_io_to_pes_4_out_valid),
    .io_to_pes_4_out_bits(PENetwork_31_io_to_pes_4_out_bits),
    .io_to_pes_5_in_valid(PENetwork_31_io_to_pes_5_in_valid),
    .io_to_pes_5_in_bits(PENetwork_31_io_to_pes_5_in_bits),
    .io_to_pes_5_out_valid(PENetwork_31_io_to_pes_5_out_valid),
    .io_to_pes_5_out_bits(PENetwork_31_io_to_pes_5_out_bits),
    .io_to_pes_6_in_valid(PENetwork_31_io_to_pes_6_in_valid),
    .io_to_pes_6_in_bits(PENetwork_31_io_to_pes_6_in_bits),
    .io_to_pes_6_out_valid(PENetwork_31_io_to_pes_6_out_valid),
    .io_to_pes_6_out_bits(PENetwork_31_io_to_pes_6_out_bits),
    .io_to_pes_7_in_valid(PENetwork_31_io_to_pes_7_in_valid),
    .io_to_pes_7_in_bits(PENetwork_31_io_to_pes_7_in_bits),
    .io_to_mem_valid(PENetwork_31_io_to_mem_valid),
    .io_to_mem_bits(PENetwork_31_io_to_mem_bits)
  );
  PENetwork_32 PENetwork_32 ( // @[pearray.scala 134:13]
    .io_to_pes_0_in_bits(PENetwork_32_io_to_pes_0_in_bits),
    .io_to_pes_0_out_bits(PENetwork_32_io_to_pes_0_out_bits),
    .io_to_pes_1_in_bits(PENetwork_32_io_to_pes_1_in_bits),
    .io_to_pes_1_out_bits(PENetwork_32_io_to_pes_1_out_bits),
    .io_to_pes_2_in_bits(PENetwork_32_io_to_pes_2_in_bits),
    .io_to_pes_2_out_bits(PENetwork_32_io_to_pes_2_out_bits),
    .io_to_pes_3_in_bits(PENetwork_32_io_to_pes_3_in_bits),
    .io_to_pes_3_out_bits(PENetwork_32_io_to_pes_3_out_bits),
    .io_to_pes_4_in_bits(PENetwork_32_io_to_pes_4_in_bits),
    .io_to_pes_4_out_bits(PENetwork_32_io_to_pes_4_out_bits),
    .io_to_pes_5_in_bits(PENetwork_32_io_to_pes_5_in_bits),
    .io_to_pes_5_out_bits(PENetwork_32_io_to_pes_5_out_bits),
    .io_to_pes_6_in_bits(PENetwork_32_io_to_pes_6_in_bits),
    .io_to_pes_6_out_bits(PENetwork_32_io_to_pes_6_out_bits),
    .io_to_pes_7_in_bits(PENetwork_32_io_to_pes_7_in_bits),
    .io_to_pes_7_out_bits(PENetwork_32_io_to_pes_7_out_bits),
    .io_to_pes_8_in_bits(PENetwork_32_io_to_pes_8_in_bits),
    .io_to_pes_8_out_bits(PENetwork_32_io_to_pes_8_out_bits),
    .io_to_pes_9_in_bits(PENetwork_32_io_to_pes_9_in_bits),
    .io_to_pes_9_out_bits(PENetwork_32_io_to_pes_9_out_bits),
    .io_to_pes_10_in_bits(PENetwork_32_io_to_pes_10_in_bits),
    .io_to_pes_10_out_bits(PENetwork_32_io_to_pes_10_out_bits),
    .io_to_pes_11_in_bits(PENetwork_32_io_to_pes_11_in_bits),
    .io_to_pes_11_out_bits(PENetwork_32_io_to_pes_11_out_bits),
    .io_to_pes_12_in_bits(PENetwork_32_io_to_pes_12_in_bits),
    .io_to_pes_12_out_bits(PENetwork_32_io_to_pes_12_out_bits),
    .io_to_pes_13_in_bits(PENetwork_32_io_to_pes_13_in_bits),
    .io_to_pes_13_out_bits(PENetwork_32_io_to_pes_13_out_bits),
    .io_to_pes_14_in_bits(PENetwork_32_io_to_pes_14_in_bits),
    .io_to_pes_14_out_bits(PENetwork_32_io_to_pes_14_out_bits),
    .io_to_pes_15_in_bits(PENetwork_32_io_to_pes_15_in_bits),
    .io_to_mem_bits(PENetwork_32_io_to_mem_bits)
  );
  PENetwork_32 PENetwork_33 ( // @[pearray.scala 134:13]
    .io_to_pes_0_in_bits(PENetwork_33_io_to_pes_0_in_bits),
    .io_to_pes_0_out_bits(PENetwork_33_io_to_pes_0_out_bits),
    .io_to_pes_1_in_bits(PENetwork_33_io_to_pes_1_in_bits),
    .io_to_pes_1_out_bits(PENetwork_33_io_to_pes_1_out_bits),
    .io_to_pes_2_in_bits(PENetwork_33_io_to_pes_2_in_bits),
    .io_to_pes_2_out_bits(PENetwork_33_io_to_pes_2_out_bits),
    .io_to_pes_3_in_bits(PENetwork_33_io_to_pes_3_in_bits),
    .io_to_pes_3_out_bits(PENetwork_33_io_to_pes_3_out_bits),
    .io_to_pes_4_in_bits(PENetwork_33_io_to_pes_4_in_bits),
    .io_to_pes_4_out_bits(PENetwork_33_io_to_pes_4_out_bits),
    .io_to_pes_5_in_bits(PENetwork_33_io_to_pes_5_in_bits),
    .io_to_pes_5_out_bits(PENetwork_33_io_to_pes_5_out_bits),
    .io_to_pes_6_in_bits(PENetwork_33_io_to_pes_6_in_bits),
    .io_to_pes_6_out_bits(PENetwork_33_io_to_pes_6_out_bits),
    .io_to_pes_7_in_bits(PENetwork_33_io_to_pes_7_in_bits),
    .io_to_pes_7_out_bits(PENetwork_33_io_to_pes_7_out_bits),
    .io_to_pes_8_in_bits(PENetwork_33_io_to_pes_8_in_bits),
    .io_to_pes_8_out_bits(PENetwork_33_io_to_pes_8_out_bits),
    .io_to_pes_9_in_bits(PENetwork_33_io_to_pes_9_in_bits),
    .io_to_pes_9_out_bits(PENetwork_33_io_to_pes_9_out_bits),
    .io_to_pes_10_in_bits(PENetwork_33_io_to_pes_10_in_bits),
    .io_to_pes_10_out_bits(PENetwork_33_io_to_pes_10_out_bits),
    .io_to_pes_11_in_bits(PENetwork_33_io_to_pes_11_in_bits),
    .io_to_pes_11_out_bits(PENetwork_33_io_to_pes_11_out_bits),
    .io_to_pes_12_in_bits(PENetwork_33_io_to_pes_12_in_bits),
    .io_to_pes_12_out_bits(PENetwork_33_io_to_pes_12_out_bits),
    .io_to_pes_13_in_bits(PENetwork_33_io_to_pes_13_in_bits),
    .io_to_pes_13_out_bits(PENetwork_33_io_to_pes_13_out_bits),
    .io_to_pes_14_in_bits(PENetwork_33_io_to_pes_14_in_bits),
    .io_to_pes_14_out_bits(PENetwork_33_io_to_pes_14_out_bits),
    .io_to_pes_15_in_bits(PENetwork_33_io_to_pes_15_in_bits),
    .io_to_mem_bits(PENetwork_33_io_to_mem_bits)
  );
  PENetwork_32 PENetwork_34 ( // @[pearray.scala 134:13]
    .io_to_pes_0_in_bits(PENetwork_34_io_to_pes_0_in_bits),
    .io_to_pes_0_out_bits(PENetwork_34_io_to_pes_0_out_bits),
    .io_to_pes_1_in_bits(PENetwork_34_io_to_pes_1_in_bits),
    .io_to_pes_1_out_bits(PENetwork_34_io_to_pes_1_out_bits),
    .io_to_pes_2_in_bits(PENetwork_34_io_to_pes_2_in_bits),
    .io_to_pes_2_out_bits(PENetwork_34_io_to_pes_2_out_bits),
    .io_to_pes_3_in_bits(PENetwork_34_io_to_pes_3_in_bits),
    .io_to_pes_3_out_bits(PENetwork_34_io_to_pes_3_out_bits),
    .io_to_pes_4_in_bits(PENetwork_34_io_to_pes_4_in_bits),
    .io_to_pes_4_out_bits(PENetwork_34_io_to_pes_4_out_bits),
    .io_to_pes_5_in_bits(PENetwork_34_io_to_pes_5_in_bits),
    .io_to_pes_5_out_bits(PENetwork_34_io_to_pes_5_out_bits),
    .io_to_pes_6_in_bits(PENetwork_34_io_to_pes_6_in_bits),
    .io_to_pes_6_out_bits(PENetwork_34_io_to_pes_6_out_bits),
    .io_to_pes_7_in_bits(PENetwork_34_io_to_pes_7_in_bits),
    .io_to_pes_7_out_bits(PENetwork_34_io_to_pes_7_out_bits),
    .io_to_pes_8_in_bits(PENetwork_34_io_to_pes_8_in_bits),
    .io_to_pes_8_out_bits(PENetwork_34_io_to_pes_8_out_bits),
    .io_to_pes_9_in_bits(PENetwork_34_io_to_pes_9_in_bits),
    .io_to_pes_9_out_bits(PENetwork_34_io_to_pes_9_out_bits),
    .io_to_pes_10_in_bits(PENetwork_34_io_to_pes_10_in_bits),
    .io_to_pes_10_out_bits(PENetwork_34_io_to_pes_10_out_bits),
    .io_to_pes_11_in_bits(PENetwork_34_io_to_pes_11_in_bits),
    .io_to_pes_11_out_bits(PENetwork_34_io_to_pes_11_out_bits),
    .io_to_pes_12_in_bits(PENetwork_34_io_to_pes_12_in_bits),
    .io_to_pes_12_out_bits(PENetwork_34_io_to_pes_12_out_bits),
    .io_to_pes_13_in_bits(PENetwork_34_io_to_pes_13_in_bits),
    .io_to_pes_13_out_bits(PENetwork_34_io_to_pes_13_out_bits),
    .io_to_pes_14_in_bits(PENetwork_34_io_to_pes_14_in_bits),
    .io_to_pes_14_out_bits(PENetwork_34_io_to_pes_14_out_bits),
    .io_to_pes_15_in_bits(PENetwork_34_io_to_pes_15_in_bits),
    .io_to_mem_bits(PENetwork_34_io_to_mem_bits)
  );
  PENetwork_32 PENetwork_35 ( // @[pearray.scala 134:13]
    .io_to_pes_0_in_bits(PENetwork_35_io_to_pes_0_in_bits),
    .io_to_pes_0_out_bits(PENetwork_35_io_to_pes_0_out_bits),
    .io_to_pes_1_in_bits(PENetwork_35_io_to_pes_1_in_bits),
    .io_to_pes_1_out_bits(PENetwork_35_io_to_pes_1_out_bits),
    .io_to_pes_2_in_bits(PENetwork_35_io_to_pes_2_in_bits),
    .io_to_pes_2_out_bits(PENetwork_35_io_to_pes_2_out_bits),
    .io_to_pes_3_in_bits(PENetwork_35_io_to_pes_3_in_bits),
    .io_to_pes_3_out_bits(PENetwork_35_io_to_pes_3_out_bits),
    .io_to_pes_4_in_bits(PENetwork_35_io_to_pes_4_in_bits),
    .io_to_pes_4_out_bits(PENetwork_35_io_to_pes_4_out_bits),
    .io_to_pes_5_in_bits(PENetwork_35_io_to_pes_5_in_bits),
    .io_to_pes_5_out_bits(PENetwork_35_io_to_pes_5_out_bits),
    .io_to_pes_6_in_bits(PENetwork_35_io_to_pes_6_in_bits),
    .io_to_pes_6_out_bits(PENetwork_35_io_to_pes_6_out_bits),
    .io_to_pes_7_in_bits(PENetwork_35_io_to_pes_7_in_bits),
    .io_to_pes_7_out_bits(PENetwork_35_io_to_pes_7_out_bits),
    .io_to_pes_8_in_bits(PENetwork_35_io_to_pes_8_in_bits),
    .io_to_pes_8_out_bits(PENetwork_35_io_to_pes_8_out_bits),
    .io_to_pes_9_in_bits(PENetwork_35_io_to_pes_9_in_bits),
    .io_to_pes_9_out_bits(PENetwork_35_io_to_pes_9_out_bits),
    .io_to_pes_10_in_bits(PENetwork_35_io_to_pes_10_in_bits),
    .io_to_pes_10_out_bits(PENetwork_35_io_to_pes_10_out_bits),
    .io_to_pes_11_in_bits(PENetwork_35_io_to_pes_11_in_bits),
    .io_to_pes_11_out_bits(PENetwork_35_io_to_pes_11_out_bits),
    .io_to_pes_12_in_bits(PENetwork_35_io_to_pes_12_in_bits),
    .io_to_pes_12_out_bits(PENetwork_35_io_to_pes_12_out_bits),
    .io_to_pes_13_in_bits(PENetwork_35_io_to_pes_13_in_bits),
    .io_to_pes_13_out_bits(PENetwork_35_io_to_pes_13_out_bits),
    .io_to_pes_14_in_bits(PENetwork_35_io_to_pes_14_in_bits),
    .io_to_pes_14_out_bits(PENetwork_35_io_to_pes_14_out_bits),
    .io_to_pes_15_in_bits(PENetwork_35_io_to_pes_15_in_bits),
    .io_to_mem_bits(PENetwork_35_io_to_mem_bits)
  );
  PENetwork_32 PENetwork_36 ( // @[pearray.scala 134:13]
    .io_to_pes_0_in_bits(PENetwork_36_io_to_pes_0_in_bits),
    .io_to_pes_0_out_bits(PENetwork_36_io_to_pes_0_out_bits),
    .io_to_pes_1_in_bits(PENetwork_36_io_to_pes_1_in_bits),
    .io_to_pes_1_out_bits(PENetwork_36_io_to_pes_1_out_bits),
    .io_to_pes_2_in_bits(PENetwork_36_io_to_pes_2_in_bits),
    .io_to_pes_2_out_bits(PENetwork_36_io_to_pes_2_out_bits),
    .io_to_pes_3_in_bits(PENetwork_36_io_to_pes_3_in_bits),
    .io_to_pes_3_out_bits(PENetwork_36_io_to_pes_3_out_bits),
    .io_to_pes_4_in_bits(PENetwork_36_io_to_pes_4_in_bits),
    .io_to_pes_4_out_bits(PENetwork_36_io_to_pes_4_out_bits),
    .io_to_pes_5_in_bits(PENetwork_36_io_to_pes_5_in_bits),
    .io_to_pes_5_out_bits(PENetwork_36_io_to_pes_5_out_bits),
    .io_to_pes_6_in_bits(PENetwork_36_io_to_pes_6_in_bits),
    .io_to_pes_6_out_bits(PENetwork_36_io_to_pes_6_out_bits),
    .io_to_pes_7_in_bits(PENetwork_36_io_to_pes_7_in_bits),
    .io_to_pes_7_out_bits(PENetwork_36_io_to_pes_7_out_bits),
    .io_to_pes_8_in_bits(PENetwork_36_io_to_pes_8_in_bits),
    .io_to_pes_8_out_bits(PENetwork_36_io_to_pes_8_out_bits),
    .io_to_pes_9_in_bits(PENetwork_36_io_to_pes_9_in_bits),
    .io_to_pes_9_out_bits(PENetwork_36_io_to_pes_9_out_bits),
    .io_to_pes_10_in_bits(PENetwork_36_io_to_pes_10_in_bits),
    .io_to_pes_10_out_bits(PENetwork_36_io_to_pes_10_out_bits),
    .io_to_pes_11_in_bits(PENetwork_36_io_to_pes_11_in_bits),
    .io_to_pes_11_out_bits(PENetwork_36_io_to_pes_11_out_bits),
    .io_to_pes_12_in_bits(PENetwork_36_io_to_pes_12_in_bits),
    .io_to_pes_12_out_bits(PENetwork_36_io_to_pes_12_out_bits),
    .io_to_pes_13_in_bits(PENetwork_36_io_to_pes_13_in_bits),
    .io_to_pes_13_out_bits(PENetwork_36_io_to_pes_13_out_bits),
    .io_to_pes_14_in_bits(PENetwork_36_io_to_pes_14_in_bits),
    .io_to_pes_14_out_bits(PENetwork_36_io_to_pes_14_out_bits),
    .io_to_pes_15_in_bits(PENetwork_36_io_to_pes_15_in_bits),
    .io_to_mem_bits(PENetwork_36_io_to_mem_bits)
  );
  PENetwork_32 PENetwork_37 ( // @[pearray.scala 134:13]
    .io_to_pes_0_in_bits(PENetwork_37_io_to_pes_0_in_bits),
    .io_to_pes_0_out_bits(PENetwork_37_io_to_pes_0_out_bits),
    .io_to_pes_1_in_bits(PENetwork_37_io_to_pes_1_in_bits),
    .io_to_pes_1_out_bits(PENetwork_37_io_to_pes_1_out_bits),
    .io_to_pes_2_in_bits(PENetwork_37_io_to_pes_2_in_bits),
    .io_to_pes_2_out_bits(PENetwork_37_io_to_pes_2_out_bits),
    .io_to_pes_3_in_bits(PENetwork_37_io_to_pes_3_in_bits),
    .io_to_pes_3_out_bits(PENetwork_37_io_to_pes_3_out_bits),
    .io_to_pes_4_in_bits(PENetwork_37_io_to_pes_4_in_bits),
    .io_to_pes_4_out_bits(PENetwork_37_io_to_pes_4_out_bits),
    .io_to_pes_5_in_bits(PENetwork_37_io_to_pes_5_in_bits),
    .io_to_pes_5_out_bits(PENetwork_37_io_to_pes_5_out_bits),
    .io_to_pes_6_in_bits(PENetwork_37_io_to_pes_6_in_bits),
    .io_to_pes_6_out_bits(PENetwork_37_io_to_pes_6_out_bits),
    .io_to_pes_7_in_bits(PENetwork_37_io_to_pes_7_in_bits),
    .io_to_pes_7_out_bits(PENetwork_37_io_to_pes_7_out_bits),
    .io_to_pes_8_in_bits(PENetwork_37_io_to_pes_8_in_bits),
    .io_to_pes_8_out_bits(PENetwork_37_io_to_pes_8_out_bits),
    .io_to_pes_9_in_bits(PENetwork_37_io_to_pes_9_in_bits),
    .io_to_pes_9_out_bits(PENetwork_37_io_to_pes_9_out_bits),
    .io_to_pes_10_in_bits(PENetwork_37_io_to_pes_10_in_bits),
    .io_to_pes_10_out_bits(PENetwork_37_io_to_pes_10_out_bits),
    .io_to_pes_11_in_bits(PENetwork_37_io_to_pes_11_in_bits),
    .io_to_pes_11_out_bits(PENetwork_37_io_to_pes_11_out_bits),
    .io_to_pes_12_in_bits(PENetwork_37_io_to_pes_12_in_bits),
    .io_to_pes_12_out_bits(PENetwork_37_io_to_pes_12_out_bits),
    .io_to_pes_13_in_bits(PENetwork_37_io_to_pes_13_in_bits),
    .io_to_pes_13_out_bits(PENetwork_37_io_to_pes_13_out_bits),
    .io_to_pes_14_in_bits(PENetwork_37_io_to_pes_14_in_bits),
    .io_to_pes_14_out_bits(PENetwork_37_io_to_pes_14_out_bits),
    .io_to_pes_15_in_bits(PENetwork_37_io_to_pes_15_in_bits),
    .io_to_mem_bits(PENetwork_37_io_to_mem_bits)
  );
  PENetwork_32 PENetwork_38 ( // @[pearray.scala 134:13]
    .io_to_pes_0_in_bits(PENetwork_38_io_to_pes_0_in_bits),
    .io_to_pes_0_out_bits(PENetwork_38_io_to_pes_0_out_bits),
    .io_to_pes_1_in_bits(PENetwork_38_io_to_pes_1_in_bits),
    .io_to_pes_1_out_bits(PENetwork_38_io_to_pes_1_out_bits),
    .io_to_pes_2_in_bits(PENetwork_38_io_to_pes_2_in_bits),
    .io_to_pes_2_out_bits(PENetwork_38_io_to_pes_2_out_bits),
    .io_to_pes_3_in_bits(PENetwork_38_io_to_pes_3_in_bits),
    .io_to_pes_3_out_bits(PENetwork_38_io_to_pes_3_out_bits),
    .io_to_pes_4_in_bits(PENetwork_38_io_to_pes_4_in_bits),
    .io_to_pes_4_out_bits(PENetwork_38_io_to_pes_4_out_bits),
    .io_to_pes_5_in_bits(PENetwork_38_io_to_pes_5_in_bits),
    .io_to_pes_5_out_bits(PENetwork_38_io_to_pes_5_out_bits),
    .io_to_pes_6_in_bits(PENetwork_38_io_to_pes_6_in_bits),
    .io_to_pes_6_out_bits(PENetwork_38_io_to_pes_6_out_bits),
    .io_to_pes_7_in_bits(PENetwork_38_io_to_pes_7_in_bits),
    .io_to_pes_7_out_bits(PENetwork_38_io_to_pes_7_out_bits),
    .io_to_pes_8_in_bits(PENetwork_38_io_to_pes_8_in_bits),
    .io_to_pes_8_out_bits(PENetwork_38_io_to_pes_8_out_bits),
    .io_to_pes_9_in_bits(PENetwork_38_io_to_pes_9_in_bits),
    .io_to_pes_9_out_bits(PENetwork_38_io_to_pes_9_out_bits),
    .io_to_pes_10_in_bits(PENetwork_38_io_to_pes_10_in_bits),
    .io_to_pes_10_out_bits(PENetwork_38_io_to_pes_10_out_bits),
    .io_to_pes_11_in_bits(PENetwork_38_io_to_pes_11_in_bits),
    .io_to_pes_11_out_bits(PENetwork_38_io_to_pes_11_out_bits),
    .io_to_pes_12_in_bits(PENetwork_38_io_to_pes_12_in_bits),
    .io_to_pes_12_out_bits(PENetwork_38_io_to_pes_12_out_bits),
    .io_to_pes_13_in_bits(PENetwork_38_io_to_pes_13_in_bits),
    .io_to_pes_13_out_bits(PENetwork_38_io_to_pes_13_out_bits),
    .io_to_pes_14_in_bits(PENetwork_38_io_to_pes_14_in_bits),
    .io_to_pes_14_out_bits(PENetwork_38_io_to_pes_14_out_bits),
    .io_to_pes_15_in_bits(PENetwork_38_io_to_pes_15_in_bits),
    .io_to_mem_bits(PENetwork_38_io_to_mem_bits)
  );
  PENetwork_32 PENetwork_39 ( // @[pearray.scala 134:13]
    .io_to_pes_0_in_bits(PENetwork_39_io_to_pes_0_in_bits),
    .io_to_pes_0_out_bits(PENetwork_39_io_to_pes_0_out_bits),
    .io_to_pes_1_in_bits(PENetwork_39_io_to_pes_1_in_bits),
    .io_to_pes_1_out_bits(PENetwork_39_io_to_pes_1_out_bits),
    .io_to_pes_2_in_bits(PENetwork_39_io_to_pes_2_in_bits),
    .io_to_pes_2_out_bits(PENetwork_39_io_to_pes_2_out_bits),
    .io_to_pes_3_in_bits(PENetwork_39_io_to_pes_3_in_bits),
    .io_to_pes_3_out_bits(PENetwork_39_io_to_pes_3_out_bits),
    .io_to_pes_4_in_bits(PENetwork_39_io_to_pes_4_in_bits),
    .io_to_pes_4_out_bits(PENetwork_39_io_to_pes_4_out_bits),
    .io_to_pes_5_in_bits(PENetwork_39_io_to_pes_5_in_bits),
    .io_to_pes_5_out_bits(PENetwork_39_io_to_pes_5_out_bits),
    .io_to_pes_6_in_bits(PENetwork_39_io_to_pes_6_in_bits),
    .io_to_pes_6_out_bits(PENetwork_39_io_to_pes_6_out_bits),
    .io_to_pes_7_in_bits(PENetwork_39_io_to_pes_7_in_bits),
    .io_to_pes_7_out_bits(PENetwork_39_io_to_pes_7_out_bits),
    .io_to_pes_8_in_bits(PENetwork_39_io_to_pes_8_in_bits),
    .io_to_pes_8_out_bits(PENetwork_39_io_to_pes_8_out_bits),
    .io_to_pes_9_in_bits(PENetwork_39_io_to_pes_9_in_bits),
    .io_to_pes_9_out_bits(PENetwork_39_io_to_pes_9_out_bits),
    .io_to_pes_10_in_bits(PENetwork_39_io_to_pes_10_in_bits),
    .io_to_pes_10_out_bits(PENetwork_39_io_to_pes_10_out_bits),
    .io_to_pes_11_in_bits(PENetwork_39_io_to_pes_11_in_bits),
    .io_to_pes_11_out_bits(PENetwork_39_io_to_pes_11_out_bits),
    .io_to_pes_12_in_bits(PENetwork_39_io_to_pes_12_in_bits),
    .io_to_pes_12_out_bits(PENetwork_39_io_to_pes_12_out_bits),
    .io_to_pes_13_in_bits(PENetwork_39_io_to_pes_13_in_bits),
    .io_to_pes_13_out_bits(PENetwork_39_io_to_pes_13_out_bits),
    .io_to_pes_14_in_bits(PENetwork_39_io_to_pes_14_in_bits),
    .io_to_pes_14_out_bits(PENetwork_39_io_to_pes_14_out_bits),
    .io_to_pes_15_in_bits(PENetwork_39_io_to_pes_15_in_bits),
    .io_to_mem_bits(PENetwork_39_io_to_mem_bits)
  );
  MemController MemController ( // @[pearray.scala 202:15]
    .clock(MemController_clock),
    .reset(MemController_reset),
    .io_rd_valid(MemController_io_rd_valid),
    .io_wr_valid(MemController_io_wr_valid),
    .io_rd_data_valid(MemController_io_rd_data_valid),
    .io_rd_data_bits(MemController_io_rd_data_bits),
    .io_wr_data_valid(MemController_io_wr_data_valid),
    .io_wr_data_bits(MemController_io_wr_data_bits)
  );
  MemController MemController_1 ( // @[pearray.scala 202:15]
    .clock(MemController_1_clock),
    .reset(MemController_1_reset),
    .io_rd_valid(MemController_1_io_rd_valid),
    .io_wr_valid(MemController_1_io_wr_valid),
    .io_rd_data_valid(MemController_1_io_rd_data_valid),
    .io_rd_data_bits(MemController_1_io_rd_data_bits),
    .io_wr_data_valid(MemController_1_io_wr_data_valid),
    .io_wr_data_bits(MemController_1_io_wr_data_bits)
  );
  MemController MemController_2 ( // @[pearray.scala 202:15]
    .clock(MemController_2_clock),
    .reset(MemController_2_reset),
    .io_rd_valid(MemController_2_io_rd_valid),
    .io_wr_valid(MemController_2_io_wr_valid),
    .io_rd_data_valid(MemController_2_io_rd_data_valid),
    .io_rd_data_bits(MemController_2_io_rd_data_bits),
    .io_wr_data_valid(MemController_2_io_wr_data_valid),
    .io_wr_data_bits(MemController_2_io_wr_data_bits)
  );
  MemController MemController_3 ( // @[pearray.scala 202:15]
    .clock(MemController_3_clock),
    .reset(MemController_3_reset),
    .io_rd_valid(MemController_3_io_rd_valid),
    .io_wr_valid(MemController_3_io_wr_valid),
    .io_rd_data_valid(MemController_3_io_rd_data_valid),
    .io_rd_data_bits(MemController_3_io_rd_data_bits),
    .io_wr_data_valid(MemController_3_io_wr_data_valid),
    .io_wr_data_bits(MemController_3_io_wr_data_bits)
  );
  MemController MemController_4 ( // @[pearray.scala 202:15]
    .clock(MemController_4_clock),
    .reset(MemController_4_reset),
    .io_rd_valid(MemController_4_io_rd_valid),
    .io_wr_valid(MemController_4_io_wr_valid),
    .io_rd_data_valid(MemController_4_io_rd_data_valid),
    .io_rd_data_bits(MemController_4_io_rd_data_bits),
    .io_wr_data_valid(MemController_4_io_wr_data_valid),
    .io_wr_data_bits(MemController_4_io_wr_data_bits)
  );
  MemController MemController_5 ( // @[pearray.scala 202:15]
    .clock(MemController_5_clock),
    .reset(MemController_5_reset),
    .io_rd_valid(MemController_5_io_rd_valid),
    .io_wr_valid(MemController_5_io_wr_valid),
    .io_rd_data_valid(MemController_5_io_rd_data_valid),
    .io_rd_data_bits(MemController_5_io_rd_data_bits),
    .io_wr_data_valid(MemController_5_io_wr_data_valid),
    .io_wr_data_bits(MemController_5_io_wr_data_bits)
  );
  MemController MemController_6 ( // @[pearray.scala 202:15]
    .clock(MemController_6_clock),
    .reset(MemController_6_reset),
    .io_rd_valid(MemController_6_io_rd_valid),
    .io_wr_valid(MemController_6_io_wr_valid),
    .io_rd_data_valid(MemController_6_io_rd_data_valid),
    .io_rd_data_bits(MemController_6_io_rd_data_bits),
    .io_wr_data_valid(MemController_6_io_wr_data_valid),
    .io_wr_data_bits(MemController_6_io_wr_data_bits)
  );
  MemController MemController_7 ( // @[pearray.scala 202:15]
    .clock(MemController_7_clock),
    .reset(MemController_7_reset),
    .io_rd_valid(MemController_7_io_rd_valid),
    .io_wr_valid(MemController_7_io_wr_valid),
    .io_rd_data_valid(MemController_7_io_rd_data_valid),
    .io_rd_data_bits(MemController_7_io_rd_data_bits),
    .io_wr_data_valid(MemController_7_io_wr_data_valid),
    .io_wr_data_bits(MemController_7_io_wr_data_bits)
  );
  MemController MemController_8 ( // @[pearray.scala 202:15]
    .clock(MemController_8_clock),
    .reset(MemController_8_reset),
    .io_rd_valid(MemController_8_io_rd_valid),
    .io_wr_valid(MemController_8_io_wr_valid),
    .io_rd_data_valid(MemController_8_io_rd_data_valid),
    .io_rd_data_bits(MemController_8_io_rd_data_bits),
    .io_wr_data_valid(MemController_8_io_wr_data_valid),
    .io_wr_data_bits(MemController_8_io_wr_data_bits)
  );
  MemController MemController_9 ( // @[pearray.scala 202:15]
    .clock(MemController_9_clock),
    .reset(MemController_9_reset),
    .io_rd_valid(MemController_9_io_rd_valid),
    .io_wr_valid(MemController_9_io_wr_valid),
    .io_rd_data_valid(MemController_9_io_rd_data_valid),
    .io_rd_data_bits(MemController_9_io_rd_data_bits),
    .io_wr_data_valid(MemController_9_io_wr_data_valid),
    .io_wr_data_bits(MemController_9_io_wr_data_bits)
  );
  MemController MemController_10 ( // @[pearray.scala 202:15]
    .clock(MemController_10_clock),
    .reset(MemController_10_reset),
    .io_rd_valid(MemController_10_io_rd_valid),
    .io_wr_valid(MemController_10_io_wr_valid),
    .io_rd_data_valid(MemController_10_io_rd_data_valid),
    .io_rd_data_bits(MemController_10_io_rd_data_bits),
    .io_wr_data_valid(MemController_10_io_wr_data_valid),
    .io_wr_data_bits(MemController_10_io_wr_data_bits)
  );
  MemController MemController_11 ( // @[pearray.scala 202:15]
    .clock(MemController_11_clock),
    .reset(MemController_11_reset),
    .io_rd_valid(MemController_11_io_rd_valid),
    .io_wr_valid(MemController_11_io_wr_valid),
    .io_rd_data_valid(MemController_11_io_rd_data_valid),
    .io_rd_data_bits(MemController_11_io_rd_data_bits),
    .io_wr_data_valid(MemController_11_io_wr_data_valid),
    .io_wr_data_bits(MemController_11_io_wr_data_bits)
  );
  MemController MemController_12 ( // @[pearray.scala 202:15]
    .clock(MemController_12_clock),
    .reset(MemController_12_reset),
    .io_rd_valid(MemController_12_io_rd_valid),
    .io_wr_valid(MemController_12_io_wr_valid),
    .io_rd_data_valid(MemController_12_io_rd_data_valid),
    .io_rd_data_bits(MemController_12_io_rd_data_bits),
    .io_wr_data_valid(MemController_12_io_wr_data_valid),
    .io_wr_data_bits(MemController_12_io_wr_data_bits)
  );
  MemController MemController_13 ( // @[pearray.scala 202:15]
    .clock(MemController_13_clock),
    .reset(MemController_13_reset),
    .io_rd_valid(MemController_13_io_rd_valid),
    .io_wr_valid(MemController_13_io_wr_valid),
    .io_rd_data_valid(MemController_13_io_rd_data_valid),
    .io_rd_data_bits(MemController_13_io_rd_data_bits),
    .io_wr_data_valid(MemController_13_io_wr_data_valid),
    .io_wr_data_bits(MemController_13_io_wr_data_bits)
  );
  MemController MemController_14 ( // @[pearray.scala 202:15]
    .clock(MemController_14_clock),
    .reset(MemController_14_reset),
    .io_rd_valid(MemController_14_io_rd_valid),
    .io_wr_valid(MemController_14_io_wr_valid),
    .io_rd_data_valid(MemController_14_io_rd_data_valid),
    .io_rd_data_bits(MemController_14_io_rd_data_bits),
    .io_wr_data_valid(MemController_14_io_wr_data_valid),
    .io_wr_data_bits(MemController_14_io_wr_data_bits)
  );
  MemController MemController_15 ( // @[pearray.scala 202:15]
    .clock(MemController_15_clock),
    .reset(MemController_15_reset),
    .io_rd_valid(MemController_15_io_rd_valid),
    .io_wr_valid(MemController_15_io_wr_valid),
    .io_rd_data_valid(MemController_15_io_rd_data_valid),
    .io_rd_data_bits(MemController_15_io_rd_data_bits),
    .io_wr_data_valid(MemController_15_io_wr_data_valid),
    .io_wr_data_bits(MemController_15_io_wr_data_bits)
  );
  MemController MemController_16 ( // @[pearray.scala 200:15]
    .clock(MemController_16_clock),
    .reset(MemController_16_reset),
    .io_rd_valid(MemController_16_io_rd_valid),
    .io_wr_valid(MemController_16_io_wr_valid),
    .io_rd_data_valid(MemController_16_io_rd_data_valid),
    .io_rd_data_bits(MemController_16_io_rd_data_bits),
    .io_wr_data_valid(MemController_16_io_wr_data_valid),
    .io_wr_data_bits(MemController_16_io_wr_data_bits)
  );
  MemController MemController_17 ( // @[pearray.scala 200:15]
    .clock(MemController_17_clock),
    .reset(MemController_17_reset),
    .io_rd_valid(MemController_17_io_rd_valid),
    .io_wr_valid(MemController_17_io_wr_valid),
    .io_rd_data_valid(MemController_17_io_rd_data_valid),
    .io_rd_data_bits(MemController_17_io_rd_data_bits),
    .io_wr_data_valid(MemController_17_io_wr_data_valid),
    .io_wr_data_bits(MemController_17_io_wr_data_bits)
  );
  MemController MemController_18 ( // @[pearray.scala 200:15]
    .clock(MemController_18_clock),
    .reset(MemController_18_reset),
    .io_rd_valid(MemController_18_io_rd_valid),
    .io_wr_valid(MemController_18_io_wr_valid),
    .io_rd_data_valid(MemController_18_io_rd_data_valid),
    .io_rd_data_bits(MemController_18_io_rd_data_bits),
    .io_wr_data_valid(MemController_18_io_wr_data_valid),
    .io_wr_data_bits(MemController_18_io_wr_data_bits)
  );
  MemController MemController_19 ( // @[pearray.scala 200:15]
    .clock(MemController_19_clock),
    .reset(MemController_19_reset),
    .io_rd_valid(MemController_19_io_rd_valid),
    .io_wr_valid(MemController_19_io_wr_valid),
    .io_rd_data_valid(MemController_19_io_rd_data_valid),
    .io_rd_data_bits(MemController_19_io_rd_data_bits),
    .io_wr_data_valid(MemController_19_io_wr_data_valid),
    .io_wr_data_bits(MemController_19_io_wr_data_bits)
  );
  MemController MemController_20 ( // @[pearray.scala 200:15]
    .clock(MemController_20_clock),
    .reset(MemController_20_reset),
    .io_rd_valid(MemController_20_io_rd_valid),
    .io_wr_valid(MemController_20_io_wr_valid),
    .io_rd_data_valid(MemController_20_io_rd_data_valid),
    .io_rd_data_bits(MemController_20_io_rd_data_bits),
    .io_wr_data_valid(MemController_20_io_wr_data_valid),
    .io_wr_data_bits(MemController_20_io_wr_data_bits)
  );
  MemController MemController_21 ( // @[pearray.scala 200:15]
    .clock(MemController_21_clock),
    .reset(MemController_21_reset),
    .io_rd_valid(MemController_21_io_rd_valid),
    .io_wr_valid(MemController_21_io_wr_valid),
    .io_rd_data_valid(MemController_21_io_rd_data_valid),
    .io_rd_data_bits(MemController_21_io_rd_data_bits),
    .io_wr_data_valid(MemController_21_io_wr_data_valid),
    .io_wr_data_bits(MemController_21_io_wr_data_bits)
  );
  MemController MemController_22 ( // @[pearray.scala 200:15]
    .clock(MemController_22_clock),
    .reset(MemController_22_reset),
    .io_rd_valid(MemController_22_io_rd_valid),
    .io_wr_valid(MemController_22_io_wr_valid),
    .io_rd_data_valid(MemController_22_io_rd_data_valid),
    .io_rd_data_bits(MemController_22_io_rd_data_bits),
    .io_wr_data_valid(MemController_22_io_wr_data_valid),
    .io_wr_data_bits(MemController_22_io_wr_data_bits)
  );
  MemController MemController_23 ( // @[pearray.scala 200:15]
    .clock(MemController_23_clock),
    .reset(MemController_23_reset),
    .io_rd_valid(MemController_23_io_rd_valid),
    .io_wr_valid(MemController_23_io_wr_valid),
    .io_rd_data_valid(MemController_23_io_rd_data_valid),
    .io_rd_data_bits(MemController_23_io_rd_data_bits),
    .io_wr_data_valid(MemController_23_io_wr_data_valid),
    .io_wr_data_bits(MemController_23_io_wr_data_bits)
  );
  MemController MemController_24 ( // @[pearray.scala 200:15]
    .clock(MemController_24_clock),
    .reset(MemController_24_reset),
    .io_rd_valid(MemController_24_io_rd_valid),
    .io_wr_valid(MemController_24_io_wr_valid),
    .io_rd_data_valid(MemController_24_io_rd_data_valid),
    .io_rd_data_bits(MemController_24_io_rd_data_bits),
    .io_wr_data_valid(MemController_24_io_wr_data_valid),
    .io_wr_data_bits(MemController_24_io_wr_data_bits)
  );
  MemController MemController_25 ( // @[pearray.scala 200:15]
    .clock(MemController_25_clock),
    .reset(MemController_25_reset),
    .io_rd_valid(MemController_25_io_rd_valid),
    .io_wr_valid(MemController_25_io_wr_valid),
    .io_rd_data_valid(MemController_25_io_rd_data_valid),
    .io_rd_data_bits(MemController_25_io_rd_data_bits),
    .io_wr_data_valid(MemController_25_io_wr_data_valid),
    .io_wr_data_bits(MemController_25_io_wr_data_bits)
  );
  MemController MemController_26 ( // @[pearray.scala 200:15]
    .clock(MemController_26_clock),
    .reset(MemController_26_reset),
    .io_rd_valid(MemController_26_io_rd_valid),
    .io_wr_valid(MemController_26_io_wr_valid),
    .io_rd_data_valid(MemController_26_io_rd_data_valid),
    .io_rd_data_bits(MemController_26_io_rd_data_bits),
    .io_wr_data_valid(MemController_26_io_wr_data_valid),
    .io_wr_data_bits(MemController_26_io_wr_data_bits)
  );
  MemController MemController_27 ( // @[pearray.scala 200:15]
    .clock(MemController_27_clock),
    .reset(MemController_27_reset),
    .io_rd_valid(MemController_27_io_rd_valid),
    .io_wr_valid(MemController_27_io_wr_valid),
    .io_rd_data_valid(MemController_27_io_rd_data_valid),
    .io_rd_data_bits(MemController_27_io_rd_data_bits),
    .io_wr_data_valid(MemController_27_io_wr_data_valid),
    .io_wr_data_bits(MemController_27_io_wr_data_bits)
  );
  MemController MemController_28 ( // @[pearray.scala 200:15]
    .clock(MemController_28_clock),
    .reset(MemController_28_reset),
    .io_rd_valid(MemController_28_io_rd_valid),
    .io_wr_valid(MemController_28_io_wr_valid),
    .io_rd_data_valid(MemController_28_io_rd_data_valid),
    .io_rd_data_bits(MemController_28_io_rd_data_bits),
    .io_wr_data_valid(MemController_28_io_wr_data_valid),
    .io_wr_data_bits(MemController_28_io_wr_data_bits)
  );
  MemController MemController_29 ( // @[pearray.scala 200:15]
    .clock(MemController_29_clock),
    .reset(MemController_29_reset),
    .io_rd_valid(MemController_29_io_rd_valid),
    .io_wr_valid(MemController_29_io_wr_valid),
    .io_rd_data_valid(MemController_29_io_rd_data_valid),
    .io_rd_data_bits(MemController_29_io_rd_data_bits),
    .io_wr_data_valid(MemController_29_io_wr_data_valid),
    .io_wr_data_bits(MemController_29_io_wr_data_bits)
  );
  MemController MemController_30 ( // @[pearray.scala 200:15]
    .clock(MemController_30_clock),
    .reset(MemController_30_reset),
    .io_rd_valid(MemController_30_io_rd_valid),
    .io_wr_valid(MemController_30_io_wr_valid),
    .io_rd_data_valid(MemController_30_io_rd_data_valid),
    .io_rd_data_bits(MemController_30_io_rd_data_bits),
    .io_wr_data_valid(MemController_30_io_wr_data_valid),
    .io_wr_data_bits(MemController_30_io_wr_data_bits)
  );
  MemController MemController_31 ( // @[pearray.scala 200:15]
    .clock(MemController_31_clock),
    .reset(MemController_31_reset),
    .io_rd_valid(MemController_31_io_rd_valid),
    .io_wr_valid(MemController_31_io_wr_valid),
    .io_rd_data_valid(MemController_31_io_rd_data_valid),
    .io_rd_data_bits(MemController_31_io_rd_data_bits),
    .io_wr_data_valid(MemController_31_io_wr_data_valid),
    .io_wr_data_bits(MemController_31_io_wr_data_bits)
  );
  MemController MemController_32 ( // @[pearray.scala 200:15]
    .clock(MemController_32_clock),
    .reset(MemController_32_reset),
    .io_rd_valid(MemController_32_io_rd_valid),
    .io_wr_valid(MemController_32_io_wr_valid),
    .io_rd_data_valid(MemController_32_io_rd_data_valid),
    .io_rd_data_bits(MemController_32_io_rd_data_bits),
    .io_wr_data_valid(MemController_32_io_wr_data_valid),
    .io_wr_data_bits(MemController_32_io_wr_data_bits)
  );
  MemController MemController_33 ( // @[pearray.scala 200:15]
    .clock(MemController_33_clock),
    .reset(MemController_33_reset),
    .io_rd_valid(MemController_33_io_rd_valid),
    .io_wr_valid(MemController_33_io_wr_valid),
    .io_rd_data_valid(MemController_33_io_rd_data_valid),
    .io_rd_data_bits(MemController_33_io_rd_data_bits),
    .io_wr_data_valid(MemController_33_io_wr_data_valid),
    .io_wr_data_bits(MemController_33_io_wr_data_bits)
  );
  MemController MemController_34 ( // @[pearray.scala 200:15]
    .clock(MemController_34_clock),
    .reset(MemController_34_reset),
    .io_rd_valid(MemController_34_io_rd_valid),
    .io_wr_valid(MemController_34_io_wr_valid),
    .io_rd_data_valid(MemController_34_io_rd_data_valid),
    .io_rd_data_bits(MemController_34_io_rd_data_bits),
    .io_wr_data_valid(MemController_34_io_wr_data_valid),
    .io_wr_data_bits(MemController_34_io_wr_data_bits)
  );
  MemController MemController_35 ( // @[pearray.scala 200:15]
    .clock(MemController_35_clock),
    .reset(MemController_35_reset),
    .io_rd_valid(MemController_35_io_rd_valid),
    .io_wr_valid(MemController_35_io_wr_valid),
    .io_rd_data_valid(MemController_35_io_rd_data_valid),
    .io_rd_data_bits(MemController_35_io_rd_data_bits),
    .io_wr_data_valid(MemController_35_io_wr_data_valid),
    .io_wr_data_bits(MemController_35_io_wr_data_bits)
  );
  MemController MemController_36 ( // @[pearray.scala 200:15]
    .clock(MemController_36_clock),
    .reset(MemController_36_reset),
    .io_rd_valid(MemController_36_io_rd_valid),
    .io_wr_valid(MemController_36_io_wr_valid),
    .io_rd_data_valid(MemController_36_io_rd_data_valid),
    .io_rd_data_bits(MemController_36_io_rd_data_bits),
    .io_wr_data_valid(MemController_36_io_wr_data_valid),
    .io_wr_data_bits(MemController_36_io_wr_data_bits)
  );
  MemController MemController_37 ( // @[pearray.scala 200:15]
    .clock(MemController_37_clock),
    .reset(MemController_37_reset),
    .io_rd_valid(MemController_37_io_rd_valid),
    .io_wr_valid(MemController_37_io_wr_valid),
    .io_rd_data_valid(MemController_37_io_rd_data_valid),
    .io_rd_data_bits(MemController_37_io_rd_data_bits),
    .io_wr_data_valid(MemController_37_io_wr_data_valid),
    .io_wr_data_bits(MemController_37_io_wr_data_bits)
  );
  MemController MemController_38 ( // @[pearray.scala 200:15]
    .clock(MemController_38_clock),
    .reset(MemController_38_reset),
    .io_rd_valid(MemController_38_io_rd_valid),
    .io_wr_valid(MemController_38_io_wr_valid),
    .io_rd_data_valid(MemController_38_io_rd_data_valid),
    .io_rd_data_bits(MemController_38_io_rd_data_bits),
    .io_wr_data_valid(MemController_38_io_wr_data_valid),
    .io_wr_data_bits(MemController_38_io_wr_data_bits)
  );
  MemController MemController_39 ( // @[pearray.scala 200:15]
    .clock(MemController_39_clock),
    .reset(MemController_39_reset),
    .io_rd_valid(MemController_39_io_rd_valid),
    .io_wr_valid(MemController_39_io_wr_valid),
    .io_rd_data_valid(MemController_39_io_rd_data_valid),
    .io_rd_data_bits(MemController_39_io_rd_data_bits),
    .io_wr_data_valid(MemController_39_io_wr_data_valid),
    .io_wr_data_bits(MemController_39_io_wr_data_bits)
  );
  assign io_data_0_out_0_valid = MemController_io_rd_data_valid; // @[pearray.scala 244:31]
  assign io_data_0_out_0_bits = MemController_io_rd_data_bits; // @[pearray.scala 244:31]
  assign io_data_0_out_1_valid = MemController_1_io_rd_data_valid; // @[pearray.scala 244:31]
  assign io_data_0_out_1_bits = MemController_1_io_rd_data_bits; // @[pearray.scala 244:31]
  assign io_data_0_out_2_valid = MemController_2_io_rd_data_valid; // @[pearray.scala 244:31]
  assign io_data_0_out_2_bits = MemController_2_io_rd_data_bits; // @[pearray.scala 244:31]
  assign io_data_0_out_3_valid = MemController_3_io_rd_data_valid; // @[pearray.scala 244:31]
  assign io_data_0_out_3_bits = MemController_3_io_rd_data_bits; // @[pearray.scala 244:31]
  assign io_data_0_out_4_valid = MemController_4_io_rd_data_valid; // @[pearray.scala 244:31]
  assign io_data_0_out_4_bits = MemController_4_io_rd_data_bits; // @[pearray.scala 244:31]
  assign io_data_0_out_5_valid = MemController_5_io_rd_data_valid; // @[pearray.scala 244:31]
  assign io_data_0_out_5_bits = MemController_5_io_rd_data_bits; // @[pearray.scala 244:31]
  assign io_data_0_out_6_valid = MemController_6_io_rd_data_valid; // @[pearray.scala 244:31]
  assign io_data_0_out_6_bits = MemController_6_io_rd_data_bits; // @[pearray.scala 244:31]
  assign io_data_0_out_7_valid = MemController_7_io_rd_data_valid; // @[pearray.scala 244:31]
  assign io_data_0_out_7_bits = MemController_7_io_rd_data_bits; // @[pearray.scala 244:31]
  assign io_data_0_out_8_valid = MemController_8_io_rd_data_valid; // @[pearray.scala 244:31]
  assign io_data_0_out_8_bits = MemController_8_io_rd_data_bits; // @[pearray.scala 244:31]
  assign io_data_0_out_9_valid = MemController_9_io_rd_data_valid; // @[pearray.scala 244:31]
  assign io_data_0_out_9_bits = MemController_9_io_rd_data_bits; // @[pearray.scala 244:31]
  assign io_data_0_out_10_valid = MemController_10_io_rd_data_valid; // @[pearray.scala 244:31]
  assign io_data_0_out_10_bits = MemController_10_io_rd_data_bits; // @[pearray.scala 244:31]
  assign io_data_0_out_11_valid = MemController_11_io_rd_data_valid; // @[pearray.scala 244:31]
  assign io_data_0_out_11_bits = MemController_11_io_rd_data_bits; // @[pearray.scala 244:31]
  assign io_data_0_out_12_valid = MemController_12_io_rd_data_valid; // @[pearray.scala 244:31]
  assign io_data_0_out_12_bits = MemController_12_io_rd_data_bits; // @[pearray.scala 244:31]
  assign io_data_0_out_13_valid = MemController_13_io_rd_data_valid; // @[pearray.scala 244:31]
  assign io_data_0_out_13_bits = MemController_13_io_rd_data_bits; // @[pearray.scala 244:31]
  assign io_data_0_out_14_valid = MemController_14_io_rd_data_valid; // @[pearray.scala 244:31]
  assign io_data_0_out_14_bits = MemController_14_io_rd_data_bits; // @[pearray.scala 244:31]
  assign io_data_0_out_15_valid = MemController_15_io_rd_data_valid; // @[pearray.scala 244:31]
  assign io_data_0_out_15_bits = MemController_15_io_rd_data_bits; // @[pearray.scala 244:31]
  assign MultiDimTime_clock = clock;
  assign MultiDimTime_reset = reset;
  assign MultiDimTime_io_in = io_exec_valid; // @[pearray.scala 146:16]
  assign PE_clock = clock;
  assign PE_reset = reset;
  assign PE_io_data_2_in_bits = PENetwork_32_io_to_pes_0_in_bits; // @[pearray.scala 157:34]
  assign PE_io_data_1_in_valid = PENetwork_16_io_to_pes_0_in_valid; // @[pearray.scala 157:34]
  assign PE_io_data_1_in_bits = PENetwork_16_io_to_pes_0_in_bits; // @[pearray.scala 157:34]
  assign PE_io_data_0_in_valid = 1'h0; // @[pearray.scala 157:34]
  assign PE_io_data_0_in_bits = 8'h0; // @[pearray.scala 157:34]
  assign PE_io_sig_stat2trans = _T_16_3; // @[pearray.scala 180:38]
  assign PE_1_clock = clock;
  assign PE_1_reset = reset;
  assign PE_1_io_data_2_in_bits = PENetwork_33_io_to_pes_0_in_bits; // @[pearray.scala 157:34]
  assign PE_1_io_data_1_in_valid = PENetwork_16_io_to_pes_1_in_valid; // @[pearray.scala 157:34]
  assign PE_1_io_data_1_in_bits = PENetwork_16_io_to_pes_1_in_bits; // @[pearray.scala 157:34]
  assign PE_1_io_data_0_in_valid = PENetwork_io_to_pes_1_in_valid; // @[pearray.scala 157:34]
  assign PE_1_io_data_0_in_bits = PENetwork_io_to_pes_1_in_bits; // @[pearray.scala 157:34]
  assign PE_1_io_sig_stat2trans = _T_28_3; // @[pearray.scala 180:38]
  assign PE_2_clock = clock;
  assign PE_2_reset = reset;
  assign PE_2_io_data_2_in_bits = PENetwork_34_io_to_pes_0_in_bits; // @[pearray.scala 157:34]
  assign PE_2_io_data_1_in_valid = PENetwork_16_io_to_pes_2_in_valid; // @[pearray.scala 157:34]
  assign PE_2_io_data_1_in_bits = PENetwork_16_io_to_pes_2_in_bits; // @[pearray.scala 157:34]
  assign PE_2_io_data_0_in_valid = PENetwork_io_to_pes_2_in_valid; // @[pearray.scala 157:34]
  assign PE_2_io_data_0_in_bits = PENetwork_io_to_pes_2_in_bits; // @[pearray.scala 157:34]
  assign PE_2_io_sig_stat2trans = _T_40_3; // @[pearray.scala 180:38]
  assign PE_3_clock = clock;
  assign PE_3_reset = reset;
  assign PE_3_io_data_2_in_bits = PENetwork_35_io_to_pes_0_in_bits; // @[pearray.scala 157:34]
  assign PE_3_io_data_1_in_valid = PENetwork_16_io_to_pes_3_in_valid; // @[pearray.scala 157:34]
  assign PE_3_io_data_1_in_bits = PENetwork_16_io_to_pes_3_in_bits; // @[pearray.scala 157:34]
  assign PE_3_io_data_0_in_valid = PENetwork_io_to_pes_3_in_valid; // @[pearray.scala 157:34]
  assign PE_3_io_data_0_in_bits = PENetwork_io_to_pes_3_in_bits; // @[pearray.scala 157:34]
  assign PE_3_io_sig_stat2trans = _T_52_3; // @[pearray.scala 180:38]
  assign PE_4_clock = clock;
  assign PE_4_reset = reset;
  assign PE_4_io_data_2_in_bits = PENetwork_36_io_to_pes_0_in_bits; // @[pearray.scala 157:34]
  assign PE_4_io_data_1_in_valid = PENetwork_16_io_to_pes_4_in_valid; // @[pearray.scala 157:34]
  assign PE_4_io_data_1_in_bits = PENetwork_16_io_to_pes_4_in_bits; // @[pearray.scala 157:34]
  assign PE_4_io_data_0_in_valid = PENetwork_io_to_pes_4_in_valid; // @[pearray.scala 157:34]
  assign PE_4_io_data_0_in_bits = PENetwork_io_to_pes_4_in_bits; // @[pearray.scala 157:34]
  assign PE_4_io_sig_stat2trans = _T_64_3; // @[pearray.scala 180:38]
  assign PE_5_clock = clock;
  assign PE_5_reset = reset;
  assign PE_5_io_data_2_in_bits = PENetwork_37_io_to_pes_0_in_bits; // @[pearray.scala 157:34]
  assign PE_5_io_data_1_in_valid = PENetwork_16_io_to_pes_5_in_valid; // @[pearray.scala 157:34]
  assign PE_5_io_data_1_in_bits = PENetwork_16_io_to_pes_5_in_bits; // @[pearray.scala 157:34]
  assign PE_5_io_data_0_in_valid = PENetwork_io_to_pes_5_in_valid; // @[pearray.scala 157:34]
  assign PE_5_io_data_0_in_bits = PENetwork_io_to_pes_5_in_bits; // @[pearray.scala 157:34]
  assign PE_5_io_sig_stat2trans = _T_76_3; // @[pearray.scala 180:38]
  assign PE_6_clock = clock;
  assign PE_6_reset = reset;
  assign PE_6_io_data_2_in_bits = PENetwork_38_io_to_pes_0_in_bits; // @[pearray.scala 157:34]
  assign PE_6_io_data_1_in_valid = PENetwork_16_io_to_pes_6_in_valid; // @[pearray.scala 157:34]
  assign PE_6_io_data_1_in_bits = PENetwork_16_io_to_pes_6_in_bits; // @[pearray.scala 157:34]
  assign PE_6_io_data_0_in_valid = PENetwork_io_to_pes_6_in_valid; // @[pearray.scala 157:34]
  assign PE_6_io_data_0_in_bits = PENetwork_io_to_pes_6_in_bits; // @[pearray.scala 157:34]
  assign PE_6_io_sig_stat2trans = _T_88_3; // @[pearray.scala 180:38]
  assign PE_7_clock = clock;
  assign PE_7_reset = reset;
  assign PE_7_io_data_2_in_bits = PENetwork_39_io_to_pes_0_in_bits; // @[pearray.scala 157:34]
  assign PE_7_io_data_1_in_valid = PENetwork_16_io_to_pes_7_in_valid; // @[pearray.scala 157:34]
  assign PE_7_io_data_1_in_bits = PENetwork_16_io_to_pes_7_in_bits; // @[pearray.scala 157:34]
  assign PE_7_io_data_0_in_valid = PENetwork_io_to_pes_7_in_valid; // @[pearray.scala 157:34]
  assign PE_7_io_data_0_in_bits = PENetwork_io_to_pes_7_in_bits; // @[pearray.scala 157:34]
  assign PE_7_io_sig_stat2trans = _T_100_3; // @[pearray.scala 180:38]
  assign PE_8_clock = clock;
  assign PE_8_reset = reset;
  assign PE_8_io_data_2_in_bits = PENetwork_32_io_to_pes_1_in_bits; // @[pearray.scala 157:34]
  assign PE_8_io_data_1_in_valid = PENetwork_17_io_to_pes_0_in_valid; // @[pearray.scala 157:34]
  assign PE_8_io_data_1_in_bits = PENetwork_17_io_to_pes_0_in_bits; // @[pearray.scala 157:34]
  assign PE_8_io_data_0_in_valid = 1'h0; // @[pearray.scala 157:34]
  assign PE_8_io_data_0_in_bits = 8'h0; // @[pearray.scala 157:34]
  assign PE_8_io_sig_stat2trans = _T_114_3; // @[pearray.scala 180:38]
  assign PE_9_clock = clock;
  assign PE_9_reset = reset;
  assign PE_9_io_data_2_in_bits = PENetwork_33_io_to_pes_1_in_bits; // @[pearray.scala 157:34]
  assign PE_9_io_data_1_in_valid = PENetwork_17_io_to_pes_1_in_valid; // @[pearray.scala 157:34]
  assign PE_9_io_data_1_in_bits = PENetwork_17_io_to_pes_1_in_bits; // @[pearray.scala 157:34]
  assign PE_9_io_data_0_in_valid = PENetwork_1_io_to_pes_1_in_valid; // @[pearray.scala 157:34]
  assign PE_9_io_data_0_in_bits = PENetwork_1_io_to_pes_1_in_bits; // @[pearray.scala 157:34]
  assign PE_9_io_sig_stat2trans = _T_126_3; // @[pearray.scala 180:38]
  assign PE_10_clock = clock;
  assign PE_10_reset = reset;
  assign PE_10_io_data_2_in_bits = PENetwork_34_io_to_pes_1_in_bits; // @[pearray.scala 157:34]
  assign PE_10_io_data_1_in_valid = PENetwork_17_io_to_pes_2_in_valid; // @[pearray.scala 157:34]
  assign PE_10_io_data_1_in_bits = PENetwork_17_io_to_pes_2_in_bits; // @[pearray.scala 157:34]
  assign PE_10_io_data_0_in_valid = PENetwork_1_io_to_pes_2_in_valid; // @[pearray.scala 157:34]
  assign PE_10_io_data_0_in_bits = PENetwork_1_io_to_pes_2_in_bits; // @[pearray.scala 157:34]
  assign PE_10_io_sig_stat2trans = _T_138_3; // @[pearray.scala 180:38]
  assign PE_11_clock = clock;
  assign PE_11_reset = reset;
  assign PE_11_io_data_2_in_bits = PENetwork_35_io_to_pes_1_in_bits; // @[pearray.scala 157:34]
  assign PE_11_io_data_1_in_valid = PENetwork_17_io_to_pes_3_in_valid; // @[pearray.scala 157:34]
  assign PE_11_io_data_1_in_bits = PENetwork_17_io_to_pes_3_in_bits; // @[pearray.scala 157:34]
  assign PE_11_io_data_0_in_valid = PENetwork_1_io_to_pes_3_in_valid; // @[pearray.scala 157:34]
  assign PE_11_io_data_0_in_bits = PENetwork_1_io_to_pes_3_in_bits; // @[pearray.scala 157:34]
  assign PE_11_io_sig_stat2trans = _T_150_3; // @[pearray.scala 180:38]
  assign PE_12_clock = clock;
  assign PE_12_reset = reset;
  assign PE_12_io_data_2_in_bits = PENetwork_36_io_to_pes_1_in_bits; // @[pearray.scala 157:34]
  assign PE_12_io_data_1_in_valid = PENetwork_17_io_to_pes_4_in_valid; // @[pearray.scala 157:34]
  assign PE_12_io_data_1_in_bits = PENetwork_17_io_to_pes_4_in_bits; // @[pearray.scala 157:34]
  assign PE_12_io_data_0_in_valid = PENetwork_1_io_to_pes_4_in_valid; // @[pearray.scala 157:34]
  assign PE_12_io_data_0_in_bits = PENetwork_1_io_to_pes_4_in_bits; // @[pearray.scala 157:34]
  assign PE_12_io_sig_stat2trans = _T_162_3; // @[pearray.scala 180:38]
  assign PE_13_clock = clock;
  assign PE_13_reset = reset;
  assign PE_13_io_data_2_in_bits = PENetwork_37_io_to_pes_1_in_bits; // @[pearray.scala 157:34]
  assign PE_13_io_data_1_in_valid = PENetwork_17_io_to_pes_5_in_valid; // @[pearray.scala 157:34]
  assign PE_13_io_data_1_in_bits = PENetwork_17_io_to_pes_5_in_bits; // @[pearray.scala 157:34]
  assign PE_13_io_data_0_in_valid = PENetwork_1_io_to_pes_5_in_valid; // @[pearray.scala 157:34]
  assign PE_13_io_data_0_in_bits = PENetwork_1_io_to_pes_5_in_bits; // @[pearray.scala 157:34]
  assign PE_13_io_sig_stat2trans = _T_174_3; // @[pearray.scala 180:38]
  assign PE_14_clock = clock;
  assign PE_14_reset = reset;
  assign PE_14_io_data_2_in_bits = PENetwork_38_io_to_pes_1_in_bits; // @[pearray.scala 157:34]
  assign PE_14_io_data_1_in_valid = PENetwork_17_io_to_pes_6_in_valid; // @[pearray.scala 157:34]
  assign PE_14_io_data_1_in_bits = PENetwork_17_io_to_pes_6_in_bits; // @[pearray.scala 157:34]
  assign PE_14_io_data_0_in_valid = PENetwork_1_io_to_pes_6_in_valid; // @[pearray.scala 157:34]
  assign PE_14_io_data_0_in_bits = PENetwork_1_io_to_pes_6_in_bits; // @[pearray.scala 157:34]
  assign PE_14_io_sig_stat2trans = _T_186_3; // @[pearray.scala 180:38]
  assign PE_15_clock = clock;
  assign PE_15_reset = reset;
  assign PE_15_io_data_2_in_bits = PENetwork_39_io_to_pes_1_in_bits; // @[pearray.scala 157:34]
  assign PE_15_io_data_1_in_valid = PENetwork_17_io_to_pes_7_in_valid; // @[pearray.scala 157:34]
  assign PE_15_io_data_1_in_bits = PENetwork_17_io_to_pes_7_in_bits; // @[pearray.scala 157:34]
  assign PE_15_io_data_0_in_valid = PENetwork_1_io_to_pes_7_in_valid; // @[pearray.scala 157:34]
  assign PE_15_io_data_0_in_bits = PENetwork_1_io_to_pes_7_in_bits; // @[pearray.scala 157:34]
  assign PE_15_io_sig_stat2trans = _T_198_3; // @[pearray.scala 180:38]
  assign PE_16_clock = clock;
  assign PE_16_reset = reset;
  assign PE_16_io_data_2_in_bits = PENetwork_32_io_to_pes_2_in_bits; // @[pearray.scala 157:34]
  assign PE_16_io_data_1_in_valid = PENetwork_18_io_to_pes_0_in_valid; // @[pearray.scala 157:34]
  assign PE_16_io_data_1_in_bits = PENetwork_18_io_to_pes_0_in_bits; // @[pearray.scala 157:34]
  assign PE_16_io_data_0_in_valid = 1'h0; // @[pearray.scala 157:34]
  assign PE_16_io_data_0_in_bits = 8'h0; // @[pearray.scala 157:34]
  assign PE_16_io_sig_stat2trans = _T_212_3; // @[pearray.scala 180:38]
  assign PE_17_clock = clock;
  assign PE_17_reset = reset;
  assign PE_17_io_data_2_in_bits = PENetwork_33_io_to_pes_2_in_bits; // @[pearray.scala 157:34]
  assign PE_17_io_data_1_in_valid = PENetwork_18_io_to_pes_1_in_valid; // @[pearray.scala 157:34]
  assign PE_17_io_data_1_in_bits = PENetwork_18_io_to_pes_1_in_bits; // @[pearray.scala 157:34]
  assign PE_17_io_data_0_in_valid = PENetwork_2_io_to_pes_1_in_valid; // @[pearray.scala 157:34]
  assign PE_17_io_data_0_in_bits = PENetwork_2_io_to_pes_1_in_bits; // @[pearray.scala 157:34]
  assign PE_17_io_sig_stat2trans = _T_224_3; // @[pearray.scala 180:38]
  assign PE_18_clock = clock;
  assign PE_18_reset = reset;
  assign PE_18_io_data_2_in_bits = PENetwork_34_io_to_pes_2_in_bits; // @[pearray.scala 157:34]
  assign PE_18_io_data_1_in_valid = PENetwork_18_io_to_pes_2_in_valid; // @[pearray.scala 157:34]
  assign PE_18_io_data_1_in_bits = PENetwork_18_io_to_pes_2_in_bits; // @[pearray.scala 157:34]
  assign PE_18_io_data_0_in_valid = PENetwork_2_io_to_pes_2_in_valid; // @[pearray.scala 157:34]
  assign PE_18_io_data_0_in_bits = PENetwork_2_io_to_pes_2_in_bits; // @[pearray.scala 157:34]
  assign PE_18_io_sig_stat2trans = _T_236_3; // @[pearray.scala 180:38]
  assign PE_19_clock = clock;
  assign PE_19_reset = reset;
  assign PE_19_io_data_2_in_bits = PENetwork_35_io_to_pes_2_in_bits; // @[pearray.scala 157:34]
  assign PE_19_io_data_1_in_valid = PENetwork_18_io_to_pes_3_in_valid; // @[pearray.scala 157:34]
  assign PE_19_io_data_1_in_bits = PENetwork_18_io_to_pes_3_in_bits; // @[pearray.scala 157:34]
  assign PE_19_io_data_0_in_valid = PENetwork_2_io_to_pes_3_in_valid; // @[pearray.scala 157:34]
  assign PE_19_io_data_0_in_bits = PENetwork_2_io_to_pes_3_in_bits; // @[pearray.scala 157:34]
  assign PE_19_io_sig_stat2trans = _T_248_3; // @[pearray.scala 180:38]
  assign PE_20_clock = clock;
  assign PE_20_reset = reset;
  assign PE_20_io_data_2_in_bits = PENetwork_36_io_to_pes_2_in_bits; // @[pearray.scala 157:34]
  assign PE_20_io_data_1_in_valid = PENetwork_18_io_to_pes_4_in_valid; // @[pearray.scala 157:34]
  assign PE_20_io_data_1_in_bits = PENetwork_18_io_to_pes_4_in_bits; // @[pearray.scala 157:34]
  assign PE_20_io_data_0_in_valid = PENetwork_2_io_to_pes_4_in_valid; // @[pearray.scala 157:34]
  assign PE_20_io_data_0_in_bits = PENetwork_2_io_to_pes_4_in_bits; // @[pearray.scala 157:34]
  assign PE_20_io_sig_stat2trans = _T_260_3; // @[pearray.scala 180:38]
  assign PE_21_clock = clock;
  assign PE_21_reset = reset;
  assign PE_21_io_data_2_in_bits = PENetwork_37_io_to_pes_2_in_bits; // @[pearray.scala 157:34]
  assign PE_21_io_data_1_in_valid = PENetwork_18_io_to_pes_5_in_valid; // @[pearray.scala 157:34]
  assign PE_21_io_data_1_in_bits = PENetwork_18_io_to_pes_5_in_bits; // @[pearray.scala 157:34]
  assign PE_21_io_data_0_in_valid = PENetwork_2_io_to_pes_5_in_valid; // @[pearray.scala 157:34]
  assign PE_21_io_data_0_in_bits = PENetwork_2_io_to_pes_5_in_bits; // @[pearray.scala 157:34]
  assign PE_21_io_sig_stat2trans = _T_272_3; // @[pearray.scala 180:38]
  assign PE_22_clock = clock;
  assign PE_22_reset = reset;
  assign PE_22_io_data_2_in_bits = PENetwork_38_io_to_pes_2_in_bits; // @[pearray.scala 157:34]
  assign PE_22_io_data_1_in_valid = PENetwork_18_io_to_pes_6_in_valid; // @[pearray.scala 157:34]
  assign PE_22_io_data_1_in_bits = PENetwork_18_io_to_pes_6_in_bits; // @[pearray.scala 157:34]
  assign PE_22_io_data_0_in_valid = PENetwork_2_io_to_pes_6_in_valid; // @[pearray.scala 157:34]
  assign PE_22_io_data_0_in_bits = PENetwork_2_io_to_pes_6_in_bits; // @[pearray.scala 157:34]
  assign PE_22_io_sig_stat2trans = _T_284_3; // @[pearray.scala 180:38]
  assign PE_23_clock = clock;
  assign PE_23_reset = reset;
  assign PE_23_io_data_2_in_bits = PENetwork_39_io_to_pes_2_in_bits; // @[pearray.scala 157:34]
  assign PE_23_io_data_1_in_valid = PENetwork_18_io_to_pes_7_in_valid; // @[pearray.scala 157:34]
  assign PE_23_io_data_1_in_bits = PENetwork_18_io_to_pes_7_in_bits; // @[pearray.scala 157:34]
  assign PE_23_io_data_0_in_valid = PENetwork_2_io_to_pes_7_in_valid; // @[pearray.scala 157:34]
  assign PE_23_io_data_0_in_bits = PENetwork_2_io_to_pes_7_in_bits; // @[pearray.scala 157:34]
  assign PE_23_io_sig_stat2trans = _T_296_3; // @[pearray.scala 180:38]
  assign PE_24_clock = clock;
  assign PE_24_reset = reset;
  assign PE_24_io_data_2_in_bits = PENetwork_32_io_to_pes_3_in_bits; // @[pearray.scala 157:34]
  assign PE_24_io_data_1_in_valid = PENetwork_19_io_to_pes_0_in_valid; // @[pearray.scala 157:34]
  assign PE_24_io_data_1_in_bits = PENetwork_19_io_to_pes_0_in_bits; // @[pearray.scala 157:34]
  assign PE_24_io_data_0_in_valid = 1'h0; // @[pearray.scala 157:34]
  assign PE_24_io_data_0_in_bits = 8'h0; // @[pearray.scala 157:34]
  assign PE_24_io_sig_stat2trans = _T_310_3; // @[pearray.scala 180:38]
  assign PE_25_clock = clock;
  assign PE_25_reset = reset;
  assign PE_25_io_data_2_in_bits = PENetwork_33_io_to_pes_3_in_bits; // @[pearray.scala 157:34]
  assign PE_25_io_data_1_in_valid = PENetwork_19_io_to_pes_1_in_valid; // @[pearray.scala 157:34]
  assign PE_25_io_data_1_in_bits = PENetwork_19_io_to_pes_1_in_bits; // @[pearray.scala 157:34]
  assign PE_25_io_data_0_in_valid = PENetwork_3_io_to_pes_1_in_valid; // @[pearray.scala 157:34]
  assign PE_25_io_data_0_in_bits = PENetwork_3_io_to_pes_1_in_bits; // @[pearray.scala 157:34]
  assign PE_25_io_sig_stat2trans = _T_322_3; // @[pearray.scala 180:38]
  assign PE_26_clock = clock;
  assign PE_26_reset = reset;
  assign PE_26_io_data_2_in_bits = PENetwork_34_io_to_pes_3_in_bits; // @[pearray.scala 157:34]
  assign PE_26_io_data_1_in_valid = PENetwork_19_io_to_pes_2_in_valid; // @[pearray.scala 157:34]
  assign PE_26_io_data_1_in_bits = PENetwork_19_io_to_pes_2_in_bits; // @[pearray.scala 157:34]
  assign PE_26_io_data_0_in_valid = PENetwork_3_io_to_pes_2_in_valid; // @[pearray.scala 157:34]
  assign PE_26_io_data_0_in_bits = PENetwork_3_io_to_pes_2_in_bits; // @[pearray.scala 157:34]
  assign PE_26_io_sig_stat2trans = _T_334_3; // @[pearray.scala 180:38]
  assign PE_27_clock = clock;
  assign PE_27_reset = reset;
  assign PE_27_io_data_2_in_bits = PENetwork_35_io_to_pes_3_in_bits; // @[pearray.scala 157:34]
  assign PE_27_io_data_1_in_valid = PENetwork_19_io_to_pes_3_in_valid; // @[pearray.scala 157:34]
  assign PE_27_io_data_1_in_bits = PENetwork_19_io_to_pes_3_in_bits; // @[pearray.scala 157:34]
  assign PE_27_io_data_0_in_valid = PENetwork_3_io_to_pes_3_in_valid; // @[pearray.scala 157:34]
  assign PE_27_io_data_0_in_bits = PENetwork_3_io_to_pes_3_in_bits; // @[pearray.scala 157:34]
  assign PE_27_io_sig_stat2trans = _T_346_3; // @[pearray.scala 180:38]
  assign PE_28_clock = clock;
  assign PE_28_reset = reset;
  assign PE_28_io_data_2_in_bits = PENetwork_36_io_to_pes_3_in_bits; // @[pearray.scala 157:34]
  assign PE_28_io_data_1_in_valid = PENetwork_19_io_to_pes_4_in_valid; // @[pearray.scala 157:34]
  assign PE_28_io_data_1_in_bits = PENetwork_19_io_to_pes_4_in_bits; // @[pearray.scala 157:34]
  assign PE_28_io_data_0_in_valid = PENetwork_3_io_to_pes_4_in_valid; // @[pearray.scala 157:34]
  assign PE_28_io_data_0_in_bits = PENetwork_3_io_to_pes_4_in_bits; // @[pearray.scala 157:34]
  assign PE_28_io_sig_stat2trans = _T_358_3; // @[pearray.scala 180:38]
  assign PE_29_clock = clock;
  assign PE_29_reset = reset;
  assign PE_29_io_data_2_in_bits = PENetwork_37_io_to_pes_3_in_bits; // @[pearray.scala 157:34]
  assign PE_29_io_data_1_in_valid = PENetwork_19_io_to_pes_5_in_valid; // @[pearray.scala 157:34]
  assign PE_29_io_data_1_in_bits = PENetwork_19_io_to_pes_5_in_bits; // @[pearray.scala 157:34]
  assign PE_29_io_data_0_in_valid = PENetwork_3_io_to_pes_5_in_valid; // @[pearray.scala 157:34]
  assign PE_29_io_data_0_in_bits = PENetwork_3_io_to_pes_5_in_bits; // @[pearray.scala 157:34]
  assign PE_29_io_sig_stat2trans = _T_370_3; // @[pearray.scala 180:38]
  assign PE_30_clock = clock;
  assign PE_30_reset = reset;
  assign PE_30_io_data_2_in_bits = PENetwork_38_io_to_pes_3_in_bits; // @[pearray.scala 157:34]
  assign PE_30_io_data_1_in_valid = PENetwork_19_io_to_pes_6_in_valid; // @[pearray.scala 157:34]
  assign PE_30_io_data_1_in_bits = PENetwork_19_io_to_pes_6_in_bits; // @[pearray.scala 157:34]
  assign PE_30_io_data_0_in_valid = PENetwork_3_io_to_pes_6_in_valid; // @[pearray.scala 157:34]
  assign PE_30_io_data_0_in_bits = PENetwork_3_io_to_pes_6_in_bits; // @[pearray.scala 157:34]
  assign PE_30_io_sig_stat2trans = _T_382_3; // @[pearray.scala 180:38]
  assign PE_31_clock = clock;
  assign PE_31_reset = reset;
  assign PE_31_io_data_2_in_bits = PENetwork_39_io_to_pes_3_in_bits; // @[pearray.scala 157:34]
  assign PE_31_io_data_1_in_valid = PENetwork_19_io_to_pes_7_in_valid; // @[pearray.scala 157:34]
  assign PE_31_io_data_1_in_bits = PENetwork_19_io_to_pes_7_in_bits; // @[pearray.scala 157:34]
  assign PE_31_io_data_0_in_valid = PENetwork_3_io_to_pes_7_in_valid; // @[pearray.scala 157:34]
  assign PE_31_io_data_0_in_bits = PENetwork_3_io_to_pes_7_in_bits; // @[pearray.scala 157:34]
  assign PE_31_io_sig_stat2trans = _T_394_3; // @[pearray.scala 180:38]
  assign PE_32_clock = clock;
  assign PE_32_reset = reset;
  assign PE_32_io_data_2_in_bits = PENetwork_32_io_to_pes_4_in_bits; // @[pearray.scala 157:34]
  assign PE_32_io_data_1_in_valid = PENetwork_20_io_to_pes_0_in_valid; // @[pearray.scala 157:34]
  assign PE_32_io_data_1_in_bits = PENetwork_20_io_to_pes_0_in_bits; // @[pearray.scala 157:34]
  assign PE_32_io_data_0_in_valid = 1'h0; // @[pearray.scala 157:34]
  assign PE_32_io_data_0_in_bits = 8'h0; // @[pearray.scala 157:34]
  assign PE_32_io_sig_stat2trans = _T_408_3; // @[pearray.scala 180:38]
  assign PE_33_clock = clock;
  assign PE_33_reset = reset;
  assign PE_33_io_data_2_in_bits = PENetwork_33_io_to_pes_4_in_bits; // @[pearray.scala 157:34]
  assign PE_33_io_data_1_in_valid = PENetwork_20_io_to_pes_1_in_valid; // @[pearray.scala 157:34]
  assign PE_33_io_data_1_in_bits = PENetwork_20_io_to_pes_1_in_bits; // @[pearray.scala 157:34]
  assign PE_33_io_data_0_in_valid = PENetwork_4_io_to_pes_1_in_valid; // @[pearray.scala 157:34]
  assign PE_33_io_data_0_in_bits = PENetwork_4_io_to_pes_1_in_bits; // @[pearray.scala 157:34]
  assign PE_33_io_sig_stat2trans = _T_420_3; // @[pearray.scala 180:38]
  assign PE_34_clock = clock;
  assign PE_34_reset = reset;
  assign PE_34_io_data_2_in_bits = PENetwork_34_io_to_pes_4_in_bits; // @[pearray.scala 157:34]
  assign PE_34_io_data_1_in_valid = PENetwork_20_io_to_pes_2_in_valid; // @[pearray.scala 157:34]
  assign PE_34_io_data_1_in_bits = PENetwork_20_io_to_pes_2_in_bits; // @[pearray.scala 157:34]
  assign PE_34_io_data_0_in_valid = PENetwork_4_io_to_pes_2_in_valid; // @[pearray.scala 157:34]
  assign PE_34_io_data_0_in_bits = PENetwork_4_io_to_pes_2_in_bits; // @[pearray.scala 157:34]
  assign PE_34_io_sig_stat2trans = _T_432_3; // @[pearray.scala 180:38]
  assign PE_35_clock = clock;
  assign PE_35_reset = reset;
  assign PE_35_io_data_2_in_bits = PENetwork_35_io_to_pes_4_in_bits; // @[pearray.scala 157:34]
  assign PE_35_io_data_1_in_valid = PENetwork_20_io_to_pes_3_in_valid; // @[pearray.scala 157:34]
  assign PE_35_io_data_1_in_bits = PENetwork_20_io_to_pes_3_in_bits; // @[pearray.scala 157:34]
  assign PE_35_io_data_0_in_valid = PENetwork_4_io_to_pes_3_in_valid; // @[pearray.scala 157:34]
  assign PE_35_io_data_0_in_bits = PENetwork_4_io_to_pes_3_in_bits; // @[pearray.scala 157:34]
  assign PE_35_io_sig_stat2trans = _T_444_3; // @[pearray.scala 180:38]
  assign PE_36_clock = clock;
  assign PE_36_reset = reset;
  assign PE_36_io_data_2_in_bits = PENetwork_36_io_to_pes_4_in_bits; // @[pearray.scala 157:34]
  assign PE_36_io_data_1_in_valid = PENetwork_20_io_to_pes_4_in_valid; // @[pearray.scala 157:34]
  assign PE_36_io_data_1_in_bits = PENetwork_20_io_to_pes_4_in_bits; // @[pearray.scala 157:34]
  assign PE_36_io_data_0_in_valid = PENetwork_4_io_to_pes_4_in_valid; // @[pearray.scala 157:34]
  assign PE_36_io_data_0_in_bits = PENetwork_4_io_to_pes_4_in_bits; // @[pearray.scala 157:34]
  assign PE_36_io_sig_stat2trans = _T_456_3; // @[pearray.scala 180:38]
  assign PE_37_clock = clock;
  assign PE_37_reset = reset;
  assign PE_37_io_data_2_in_bits = PENetwork_37_io_to_pes_4_in_bits; // @[pearray.scala 157:34]
  assign PE_37_io_data_1_in_valid = PENetwork_20_io_to_pes_5_in_valid; // @[pearray.scala 157:34]
  assign PE_37_io_data_1_in_bits = PENetwork_20_io_to_pes_5_in_bits; // @[pearray.scala 157:34]
  assign PE_37_io_data_0_in_valid = PENetwork_4_io_to_pes_5_in_valid; // @[pearray.scala 157:34]
  assign PE_37_io_data_0_in_bits = PENetwork_4_io_to_pes_5_in_bits; // @[pearray.scala 157:34]
  assign PE_37_io_sig_stat2trans = _T_468_3; // @[pearray.scala 180:38]
  assign PE_38_clock = clock;
  assign PE_38_reset = reset;
  assign PE_38_io_data_2_in_bits = PENetwork_38_io_to_pes_4_in_bits; // @[pearray.scala 157:34]
  assign PE_38_io_data_1_in_valid = PENetwork_20_io_to_pes_6_in_valid; // @[pearray.scala 157:34]
  assign PE_38_io_data_1_in_bits = PENetwork_20_io_to_pes_6_in_bits; // @[pearray.scala 157:34]
  assign PE_38_io_data_0_in_valid = PENetwork_4_io_to_pes_6_in_valid; // @[pearray.scala 157:34]
  assign PE_38_io_data_0_in_bits = PENetwork_4_io_to_pes_6_in_bits; // @[pearray.scala 157:34]
  assign PE_38_io_sig_stat2trans = _T_480_3; // @[pearray.scala 180:38]
  assign PE_39_clock = clock;
  assign PE_39_reset = reset;
  assign PE_39_io_data_2_in_bits = PENetwork_39_io_to_pes_4_in_bits; // @[pearray.scala 157:34]
  assign PE_39_io_data_1_in_valid = PENetwork_20_io_to_pes_7_in_valid; // @[pearray.scala 157:34]
  assign PE_39_io_data_1_in_bits = PENetwork_20_io_to_pes_7_in_bits; // @[pearray.scala 157:34]
  assign PE_39_io_data_0_in_valid = PENetwork_4_io_to_pes_7_in_valid; // @[pearray.scala 157:34]
  assign PE_39_io_data_0_in_bits = PENetwork_4_io_to_pes_7_in_bits; // @[pearray.scala 157:34]
  assign PE_39_io_sig_stat2trans = _T_492_3; // @[pearray.scala 180:38]
  assign PE_40_clock = clock;
  assign PE_40_reset = reset;
  assign PE_40_io_data_2_in_bits = PENetwork_32_io_to_pes_5_in_bits; // @[pearray.scala 157:34]
  assign PE_40_io_data_1_in_valid = PENetwork_21_io_to_pes_0_in_valid; // @[pearray.scala 157:34]
  assign PE_40_io_data_1_in_bits = PENetwork_21_io_to_pes_0_in_bits; // @[pearray.scala 157:34]
  assign PE_40_io_data_0_in_valid = 1'h0; // @[pearray.scala 157:34]
  assign PE_40_io_data_0_in_bits = 8'h0; // @[pearray.scala 157:34]
  assign PE_40_io_sig_stat2trans = _T_506_3; // @[pearray.scala 180:38]
  assign PE_41_clock = clock;
  assign PE_41_reset = reset;
  assign PE_41_io_data_2_in_bits = PENetwork_33_io_to_pes_5_in_bits; // @[pearray.scala 157:34]
  assign PE_41_io_data_1_in_valid = PENetwork_21_io_to_pes_1_in_valid; // @[pearray.scala 157:34]
  assign PE_41_io_data_1_in_bits = PENetwork_21_io_to_pes_1_in_bits; // @[pearray.scala 157:34]
  assign PE_41_io_data_0_in_valid = PENetwork_5_io_to_pes_1_in_valid; // @[pearray.scala 157:34]
  assign PE_41_io_data_0_in_bits = PENetwork_5_io_to_pes_1_in_bits; // @[pearray.scala 157:34]
  assign PE_41_io_sig_stat2trans = _T_518_3; // @[pearray.scala 180:38]
  assign PE_42_clock = clock;
  assign PE_42_reset = reset;
  assign PE_42_io_data_2_in_bits = PENetwork_34_io_to_pes_5_in_bits; // @[pearray.scala 157:34]
  assign PE_42_io_data_1_in_valid = PENetwork_21_io_to_pes_2_in_valid; // @[pearray.scala 157:34]
  assign PE_42_io_data_1_in_bits = PENetwork_21_io_to_pes_2_in_bits; // @[pearray.scala 157:34]
  assign PE_42_io_data_0_in_valid = PENetwork_5_io_to_pes_2_in_valid; // @[pearray.scala 157:34]
  assign PE_42_io_data_0_in_bits = PENetwork_5_io_to_pes_2_in_bits; // @[pearray.scala 157:34]
  assign PE_42_io_sig_stat2trans = _T_530_3; // @[pearray.scala 180:38]
  assign PE_43_clock = clock;
  assign PE_43_reset = reset;
  assign PE_43_io_data_2_in_bits = PENetwork_35_io_to_pes_5_in_bits; // @[pearray.scala 157:34]
  assign PE_43_io_data_1_in_valid = PENetwork_21_io_to_pes_3_in_valid; // @[pearray.scala 157:34]
  assign PE_43_io_data_1_in_bits = PENetwork_21_io_to_pes_3_in_bits; // @[pearray.scala 157:34]
  assign PE_43_io_data_0_in_valid = PENetwork_5_io_to_pes_3_in_valid; // @[pearray.scala 157:34]
  assign PE_43_io_data_0_in_bits = PENetwork_5_io_to_pes_3_in_bits; // @[pearray.scala 157:34]
  assign PE_43_io_sig_stat2trans = _T_542_3; // @[pearray.scala 180:38]
  assign PE_44_clock = clock;
  assign PE_44_reset = reset;
  assign PE_44_io_data_2_in_bits = PENetwork_36_io_to_pes_5_in_bits; // @[pearray.scala 157:34]
  assign PE_44_io_data_1_in_valid = PENetwork_21_io_to_pes_4_in_valid; // @[pearray.scala 157:34]
  assign PE_44_io_data_1_in_bits = PENetwork_21_io_to_pes_4_in_bits; // @[pearray.scala 157:34]
  assign PE_44_io_data_0_in_valid = PENetwork_5_io_to_pes_4_in_valid; // @[pearray.scala 157:34]
  assign PE_44_io_data_0_in_bits = PENetwork_5_io_to_pes_4_in_bits; // @[pearray.scala 157:34]
  assign PE_44_io_sig_stat2trans = _T_554_3; // @[pearray.scala 180:38]
  assign PE_45_clock = clock;
  assign PE_45_reset = reset;
  assign PE_45_io_data_2_in_bits = PENetwork_37_io_to_pes_5_in_bits; // @[pearray.scala 157:34]
  assign PE_45_io_data_1_in_valid = PENetwork_21_io_to_pes_5_in_valid; // @[pearray.scala 157:34]
  assign PE_45_io_data_1_in_bits = PENetwork_21_io_to_pes_5_in_bits; // @[pearray.scala 157:34]
  assign PE_45_io_data_0_in_valid = PENetwork_5_io_to_pes_5_in_valid; // @[pearray.scala 157:34]
  assign PE_45_io_data_0_in_bits = PENetwork_5_io_to_pes_5_in_bits; // @[pearray.scala 157:34]
  assign PE_45_io_sig_stat2trans = _T_566_3; // @[pearray.scala 180:38]
  assign PE_46_clock = clock;
  assign PE_46_reset = reset;
  assign PE_46_io_data_2_in_bits = PENetwork_38_io_to_pes_5_in_bits; // @[pearray.scala 157:34]
  assign PE_46_io_data_1_in_valid = PENetwork_21_io_to_pes_6_in_valid; // @[pearray.scala 157:34]
  assign PE_46_io_data_1_in_bits = PENetwork_21_io_to_pes_6_in_bits; // @[pearray.scala 157:34]
  assign PE_46_io_data_0_in_valid = PENetwork_5_io_to_pes_6_in_valid; // @[pearray.scala 157:34]
  assign PE_46_io_data_0_in_bits = PENetwork_5_io_to_pes_6_in_bits; // @[pearray.scala 157:34]
  assign PE_46_io_sig_stat2trans = _T_578_3; // @[pearray.scala 180:38]
  assign PE_47_clock = clock;
  assign PE_47_reset = reset;
  assign PE_47_io_data_2_in_bits = PENetwork_39_io_to_pes_5_in_bits; // @[pearray.scala 157:34]
  assign PE_47_io_data_1_in_valid = PENetwork_21_io_to_pes_7_in_valid; // @[pearray.scala 157:34]
  assign PE_47_io_data_1_in_bits = PENetwork_21_io_to_pes_7_in_bits; // @[pearray.scala 157:34]
  assign PE_47_io_data_0_in_valid = PENetwork_5_io_to_pes_7_in_valid; // @[pearray.scala 157:34]
  assign PE_47_io_data_0_in_bits = PENetwork_5_io_to_pes_7_in_bits; // @[pearray.scala 157:34]
  assign PE_47_io_sig_stat2trans = _T_590_3; // @[pearray.scala 180:38]
  assign PE_48_clock = clock;
  assign PE_48_reset = reset;
  assign PE_48_io_data_2_in_bits = PENetwork_32_io_to_pes_6_in_bits; // @[pearray.scala 157:34]
  assign PE_48_io_data_1_in_valid = PENetwork_22_io_to_pes_0_in_valid; // @[pearray.scala 157:34]
  assign PE_48_io_data_1_in_bits = PENetwork_22_io_to_pes_0_in_bits; // @[pearray.scala 157:34]
  assign PE_48_io_data_0_in_valid = 1'h0; // @[pearray.scala 157:34]
  assign PE_48_io_data_0_in_bits = 8'h0; // @[pearray.scala 157:34]
  assign PE_48_io_sig_stat2trans = _T_604_3; // @[pearray.scala 180:38]
  assign PE_49_clock = clock;
  assign PE_49_reset = reset;
  assign PE_49_io_data_2_in_bits = PENetwork_33_io_to_pes_6_in_bits; // @[pearray.scala 157:34]
  assign PE_49_io_data_1_in_valid = PENetwork_22_io_to_pes_1_in_valid; // @[pearray.scala 157:34]
  assign PE_49_io_data_1_in_bits = PENetwork_22_io_to_pes_1_in_bits; // @[pearray.scala 157:34]
  assign PE_49_io_data_0_in_valid = PENetwork_6_io_to_pes_1_in_valid; // @[pearray.scala 157:34]
  assign PE_49_io_data_0_in_bits = PENetwork_6_io_to_pes_1_in_bits; // @[pearray.scala 157:34]
  assign PE_49_io_sig_stat2trans = _T_616_3; // @[pearray.scala 180:38]
  assign PE_50_clock = clock;
  assign PE_50_reset = reset;
  assign PE_50_io_data_2_in_bits = PENetwork_34_io_to_pes_6_in_bits; // @[pearray.scala 157:34]
  assign PE_50_io_data_1_in_valid = PENetwork_22_io_to_pes_2_in_valid; // @[pearray.scala 157:34]
  assign PE_50_io_data_1_in_bits = PENetwork_22_io_to_pes_2_in_bits; // @[pearray.scala 157:34]
  assign PE_50_io_data_0_in_valid = PENetwork_6_io_to_pes_2_in_valid; // @[pearray.scala 157:34]
  assign PE_50_io_data_0_in_bits = PENetwork_6_io_to_pes_2_in_bits; // @[pearray.scala 157:34]
  assign PE_50_io_sig_stat2trans = _T_628_3; // @[pearray.scala 180:38]
  assign PE_51_clock = clock;
  assign PE_51_reset = reset;
  assign PE_51_io_data_2_in_bits = PENetwork_35_io_to_pes_6_in_bits; // @[pearray.scala 157:34]
  assign PE_51_io_data_1_in_valid = PENetwork_22_io_to_pes_3_in_valid; // @[pearray.scala 157:34]
  assign PE_51_io_data_1_in_bits = PENetwork_22_io_to_pes_3_in_bits; // @[pearray.scala 157:34]
  assign PE_51_io_data_0_in_valid = PENetwork_6_io_to_pes_3_in_valid; // @[pearray.scala 157:34]
  assign PE_51_io_data_0_in_bits = PENetwork_6_io_to_pes_3_in_bits; // @[pearray.scala 157:34]
  assign PE_51_io_sig_stat2trans = _T_640_3; // @[pearray.scala 180:38]
  assign PE_52_clock = clock;
  assign PE_52_reset = reset;
  assign PE_52_io_data_2_in_bits = PENetwork_36_io_to_pes_6_in_bits; // @[pearray.scala 157:34]
  assign PE_52_io_data_1_in_valid = PENetwork_22_io_to_pes_4_in_valid; // @[pearray.scala 157:34]
  assign PE_52_io_data_1_in_bits = PENetwork_22_io_to_pes_4_in_bits; // @[pearray.scala 157:34]
  assign PE_52_io_data_0_in_valid = PENetwork_6_io_to_pes_4_in_valid; // @[pearray.scala 157:34]
  assign PE_52_io_data_0_in_bits = PENetwork_6_io_to_pes_4_in_bits; // @[pearray.scala 157:34]
  assign PE_52_io_sig_stat2trans = _T_652_3; // @[pearray.scala 180:38]
  assign PE_53_clock = clock;
  assign PE_53_reset = reset;
  assign PE_53_io_data_2_in_bits = PENetwork_37_io_to_pes_6_in_bits; // @[pearray.scala 157:34]
  assign PE_53_io_data_1_in_valid = PENetwork_22_io_to_pes_5_in_valid; // @[pearray.scala 157:34]
  assign PE_53_io_data_1_in_bits = PENetwork_22_io_to_pes_5_in_bits; // @[pearray.scala 157:34]
  assign PE_53_io_data_0_in_valid = PENetwork_6_io_to_pes_5_in_valid; // @[pearray.scala 157:34]
  assign PE_53_io_data_0_in_bits = PENetwork_6_io_to_pes_5_in_bits; // @[pearray.scala 157:34]
  assign PE_53_io_sig_stat2trans = _T_664_3; // @[pearray.scala 180:38]
  assign PE_54_clock = clock;
  assign PE_54_reset = reset;
  assign PE_54_io_data_2_in_bits = PENetwork_38_io_to_pes_6_in_bits; // @[pearray.scala 157:34]
  assign PE_54_io_data_1_in_valid = PENetwork_22_io_to_pes_6_in_valid; // @[pearray.scala 157:34]
  assign PE_54_io_data_1_in_bits = PENetwork_22_io_to_pes_6_in_bits; // @[pearray.scala 157:34]
  assign PE_54_io_data_0_in_valid = PENetwork_6_io_to_pes_6_in_valid; // @[pearray.scala 157:34]
  assign PE_54_io_data_0_in_bits = PENetwork_6_io_to_pes_6_in_bits; // @[pearray.scala 157:34]
  assign PE_54_io_sig_stat2trans = _T_676_3; // @[pearray.scala 180:38]
  assign PE_55_clock = clock;
  assign PE_55_reset = reset;
  assign PE_55_io_data_2_in_bits = PENetwork_39_io_to_pes_6_in_bits; // @[pearray.scala 157:34]
  assign PE_55_io_data_1_in_valid = PENetwork_22_io_to_pes_7_in_valid; // @[pearray.scala 157:34]
  assign PE_55_io_data_1_in_bits = PENetwork_22_io_to_pes_7_in_bits; // @[pearray.scala 157:34]
  assign PE_55_io_data_0_in_valid = PENetwork_6_io_to_pes_7_in_valid; // @[pearray.scala 157:34]
  assign PE_55_io_data_0_in_bits = PENetwork_6_io_to_pes_7_in_bits; // @[pearray.scala 157:34]
  assign PE_55_io_sig_stat2trans = _T_688_3; // @[pearray.scala 180:38]
  assign PE_56_clock = clock;
  assign PE_56_reset = reset;
  assign PE_56_io_data_2_in_bits = PENetwork_32_io_to_pes_7_in_bits; // @[pearray.scala 157:34]
  assign PE_56_io_data_1_in_valid = PENetwork_23_io_to_pes_0_in_valid; // @[pearray.scala 157:34]
  assign PE_56_io_data_1_in_bits = PENetwork_23_io_to_pes_0_in_bits; // @[pearray.scala 157:34]
  assign PE_56_io_data_0_in_valid = 1'h0; // @[pearray.scala 157:34]
  assign PE_56_io_data_0_in_bits = 8'h0; // @[pearray.scala 157:34]
  assign PE_56_io_sig_stat2trans = _T_702_3; // @[pearray.scala 180:38]
  assign PE_57_clock = clock;
  assign PE_57_reset = reset;
  assign PE_57_io_data_2_in_bits = PENetwork_33_io_to_pes_7_in_bits; // @[pearray.scala 157:34]
  assign PE_57_io_data_1_in_valid = PENetwork_23_io_to_pes_1_in_valid; // @[pearray.scala 157:34]
  assign PE_57_io_data_1_in_bits = PENetwork_23_io_to_pes_1_in_bits; // @[pearray.scala 157:34]
  assign PE_57_io_data_0_in_valid = PENetwork_7_io_to_pes_1_in_valid; // @[pearray.scala 157:34]
  assign PE_57_io_data_0_in_bits = PENetwork_7_io_to_pes_1_in_bits; // @[pearray.scala 157:34]
  assign PE_57_io_sig_stat2trans = _T_714_3; // @[pearray.scala 180:38]
  assign PE_58_clock = clock;
  assign PE_58_reset = reset;
  assign PE_58_io_data_2_in_bits = PENetwork_34_io_to_pes_7_in_bits; // @[pearray.scala 157:34]
  assign PE_58_io_data_1_in_valid = PENetwork_23_io_to_pes_2_in_valid; // @[pearray.scala 157:34]
  assign PE_58_io_data_1_in_bits = PENetwork_23_io_to_pes_2_in_bits; // @[pearray.scala 157:34]
  assign PE_58_io_data_0_in_valid = PENetwork_7_io_to_pes_2_in_valid; // @[pearray.scala 157:34]
  assign PE_58_io_data_0_in_bits = PENetwork_7_io_to_pes_2_in_bits; // @[pearray.scala 157:34]
  assign PE_58_io_sig_stat2trans = _T_726_3; // @[pearray.scala 180:38]
  assign PE_59_clock = clock;
  assign PE_59_reset = reset;
  assign PE_59_io_data_2_in_bits = PENetwork_35_io_to_pes_7_in_bits; // @[pearray.scala 157:34]
  assign PE_59_io_data_1_in_valid = PENetwork_23_io_to_pes_3_in_valid; // @[pearray.scala 157:34]
  assign PE_59_io_data_1_in_bits = PENetwork_23_io_to_pes_3_in_bits; // @[pearray.scala 157:34]
  assign PE_59_io_data_0_in_valid = PENetwork_7_io_to_pes_3_in_valid; // @[pearray.scala 157:34]
  assign PE_59_io_data_0_in_bits = PENetwork_7_io_to_pes_3_in_bits; // @[pearray.scala 157:34]
  assign PE_59_io_sig_stat2trans = _T_738_3; // @[pearray.scala 180:38]
  assign PE_60_clock = clock;
  assign PE_60_reset = reset;
  assign PE_60_io_data_2_in_bits = PENetwork_36_io_to_pes_7_in_bits; // @[pearray.scala 157:34]
  assign PE_60_io_data_1_in_valid = PENetwork_23_io_to_pes_4_in_valid; // @[pearray.scala 157:34]
  assign PE_60_io_data_1_in_bits = PENetwork_23_io_to_pes_4_in_bits; // @[pearray.scala 157:34]
  assign PE_60_io_data_0_in_valid = PENetwork_7_io_to_pes_4_in_valid; // @[pearray.scala 157:34]
  assign PE_60_io_data_0_in_bits = PENetwork_7_io_to_pes_4_in_bits; // @[pearray.scala 157:34]
  assign PE_60_io_sig_stat2trans = _T_750_3; // @[pearray.scala 180:38]
  assign PE_61_clock = clock;
  assign PE_61_reset = reset;
  assign PE_61_io_data_2_in_bits = PENetwork_37_io_to_pes_7_in_bits; // @[pearray.scala 157:34]
  assign PE_61_io_data_1_in_valid = PENetwork_23_io_to_pes_5_in_valid; // @[pearray.scala 157:34]
  assign PE_61_io_data_1_in_bits = PENetwork_23_io_to_pes_5_in_bits; // @[pearray.scala 157:34]
  assign PE_61_io_data_0_in_valid = PENetwork_7_io_to_pes_5_in_valid; // @[pearray.scala 157:34]
  assign PE_61_io_data_0_in_bits = PENetwork_7_io_to_pes_5_in_bits; // @[pearray.scala 157:34]
  assign PE_61_io_sig_stat2trans = _T_762_3; // @[pearray.scala 180:38]
  assign PE_62_clock = clock;
  assign PE_62_reset = reset;
  assign PE_62_io_data_2_in_bits = PENetwork_38_io_to_pes_7_in_bits; // @[pearray.scala 157:34]
  assign PE_62_io_data_1_in_valid = PENetwork_23_io_to_pes_6_in_valid; // @[pearray.scala 157:34]
  assign PE_62_io_data_1_in_bits = PENetwork_23_io_to_pes_6_in_bits; // @[pearray.scala 157:34]
  assign PE_62_io_data_0_in_valid = PENetwork_7_io_to_pes_6_in_valid; // @[pearray.scala 157:34]
  assign PE_62_io_data_0_in_bits = PENetwork_7_io_to_pes_6_in_bits; // @[pearray.scala 157:34]
  assign PE_62_io_sig_stat2trans = _T_774_3; // @[pearray.scala 180:38]
  assign PE_63_clock = clock;
  assign PE_63_reset = reset;
  assign PE_63_io_data_2_in_bits = PENetwork_39_io_to_pes_7_in_bits; // @[pearray.scala 157:34]
  assign PE_63_io_data_1_in_valid = PENetwork_23_io_to_pes_7_in_valid; // @[pearray.scala 157:34]
  assign PE_63_io_data_1_in_bits = PENetwork_23_io_to_pes_7_in_bits; // @[pearray.scala 157:34]
  assign PE_63_io_data_0_in_valid = PENetwork_7_io_to_pes_7_in_valid; // @[pearray.scala 157:34]
  assign PE_63_io_data_0_in_bits = PENetwork_7_io_to_pes_7_in_bits; // @[pearray.scala 157:34]
  assign PE_63_io_sig_stat2trans = _T_786_3; // @[pearray.scala 180:38]
  assign PE_64_clock = clock;
  assign PE_64_reset = reset;
  assign PE_64_io_data_2_in_bits = PENetwork_32_io_to_pes_8_in_bits; // @[pearray.scala 157:34]
  assign PE_64_io_data_1_in_valid = PENetwork_24_io_to_pes_0_in_valid; // @[pearray.scala 157:34]
  assign PE_64_io_data_1_in_bits = PENetwork_24_io_to_pes_0_in_bits; // @[pearray.scala 157:34]
  assign PE_64_io_data_0_in_valid = 1'h0; // @[pearray.scala 157:34]
  assign PE_64_io_data_0_in_bits = 8'h0; // @[pearray.scala 157:34]
  assign PE_64_io_sig_stat2trans = _T_800_3; // @[pearray.scala 180:38]
  assign PE_65_clock = clock;
  assign PE_65_reset = reset;
  assign PE_65_io_data_2_in_bits = PENetwork_33_io_to_pes_8_in_bits; // @[pearray.scala 157:34]
  assign PE_65_io_data_1_in_valid = PENetwork_24_io_to_pes_1_in_valid; // @[pearray.scala 157:34]
  assign PE_65_io_data_1_in_bits = PENetwork_24_io_to_pes_1_in_bits; // @[pearray.scala 157:34]
  assign PE_65_io_data_0_in_valid = PENetwork_8_io_to_pes_1_in_valid; // @[pearray.scala 157:34]
  assign PE_65_io_data_0_in_bits = PENetwork_8_io_to_pes_1_in_bits; // @[pearray.scala 157:34]
  assign PE_65_io_sig_stat2trans = _T_812_3; // @[pearray.scala 180:38]
  assign PE_66_clock = clock;
  assign PE_66_reset = reset;
  assign PE_66_io_data_2_in_bits = PENetwork_34_io_to_pes_8_in_bits; // @[pearray.scala 157:34]
  assign PE_66_io_data_1_in_valid = PENetwork_24_io_to_pes_2_in_valid; // @[pearray.scala 157:34]
  assign PE_66_io_data_1_in_bits = PENetwork_24_io_to_pes_2_in_bits; // @[pearray.scala 157:34]
  assign PE_66_io_data_0_in_valid = PENetwork_8_io_to_pes_2_in_valid; // @[pearray.scala 157:34]
  assign PE_66_io_data_0_in_bits = PENetwork_8_io_to_pes_2_in_bits; // @[pearray.scala 157:34]
  assign PE_66_io_sig_stat2trans = _T_824_3; // @[pearray.scala 180:38]
  assign PE_67_clock = clock;
  assign PE_67_reset = reset;
  assign PE_67_io_data_2_in_bits = PENetwork_35_io_to_pes_8_in_bits; // @[pearray.scala 157:34]
  assign PE_67_io_data_1_in_valid = PENetwork_24_io_to_pes_3_in_valid; // @[pearray.scala 157:34]
  assign PE_67_io_data_1_in_bits = PENetwork_24_io_to_pes_3_in_bits; // @[pearray.scala 157:34]
  assign PE_67_io_data_0_in_valid = PENetwork_8_io_to_pes_3_in_valid; // @[pearray.scala 157:34]
  assign PE_67_io_data_0_in_bits = PENetwork_8_io_to_pes_3_in_bits; // @[pearray.scala 157:34]
  assign PE_67_io_sig_stat2trans = _T_836_3; // @[pearray.scala 180:38]
  assign PE_68_clock = clock;
  assign PE_68_reset = reset;
  assign PE_68_io_data_2_in_bits = PENetwork_36_io_to_pes_8_in_bits; // @[pearray.scala 157:34]
  assign PE_68_io_data_1_in_valid = PENetwork_24_io_to_pes_4_in_valid; // @[pearray.scala 157:34]
  assign PE_68_io_data_1_in_bits = PENetwork_24_io_to_pes_4_in_bits; // @[pearray.scala 157:34]
  assign PE_68_io_data_0_in_valid = PENetwork_8_io_to_pes_4_in_valid; // @[pearray.scala 157:34]
  assign PE_68_io_data_0_in_bits = PENetwork_8_io_to_pes_4_in_bits; // @[pearray.scala 157:34]
  assign PE_68_io_sig_stat2trans = _T_848_3; // @[pearray.scala 180:38]
  assign PE_69_clock = clock;
  assign PE_69_reset = reset;
  assign PE_69_io_data_2_in_bits = PENetwork_37_io_to_pes_8_in_bits; // @[pearray.scala 157:34]
  assign PE_69_io_data_1_in_valid = PENetwork_24_io_to_pes_5_in_valid; // @[pearray.scala 157:34]
  assign PE_69_io_data_1_in_bits = PENetwork_24_io_to_pes_5_in_bits; // @[pearray.scala 157:34]
  assign PE_69_io_data_0_in_valid = PENetwork_8_io_to_pes_5_in_valid; // @[pearray.scala 157:34]
  assign PE_69_io_data_0_in_bits = PENetwork_8_io_to_pes_5_in_bits; // @[pearray.scala 157:34]
  assign PE_69_io_sig_stat2trans = _T_860_3; // @[pearray.scala 180:38]
  assign PE_70_clock = clock;
  assign PE_70_reset = reset;
  assign PE_70_io_data_2_in_bits = PENetwork_38_io_to_pes_8_in_bits; // @[pearray.scala 157:34]
  assign PE_70_io_data_1_in_valid = PENetwork_24_io_to_pes_6_in_valid; // @[pearray.scala 157:34]
  assign PE_70_io_data_1_in_bits = PENetwork_24_io_to_pes_6_in_bits; // @[pearray.scala 157:34]
  assign PE_70_io_data_0_in_valid = PENetwork_8_io_to_pes_6_in_valid; // @[pearray.scala 157:34]
  assign PE_70_io_data_0_in_bits = PENetwork_8_io_to_pes_6_in_bits; // @[pearray.scala 157:34]
  assign PE_70_io_sig_stat2trans = _T_872_3; // @[pearray.scala 180:38]
  assign PE_71_clock = clock;
  assign PE_71_reset = reset;
  assign PE_71_io_data_2_in_bits = PENetwork_39_io_to_pes_8_in_bits; // @[pearray.scala 157:34]
  assign PE_71_io_data_1_in_valid = PENetwork_24_io_to_pes_7_in_valid; // @[pearray.scala 157:34]
  assign PE_71_io_data_1_in_bits = PENetwork_24_io_to_pes_7_in_bits; // @[pearray.scala 157:34]
  assign PE_71_io_data_0_in_valid = PENetwork_8_io_to_pes_7_in_valid; // @[pearray.scala 157:34]
  assign PE_71_io_data_0_in_bits = PENetwork_8_io_to_pes_7_in_bits; // @[pearray.scala 157:34]
  assign PE_71_io_sig_stat2trans = _T_884_3; // @[pearray.scala 180:38]
  assign PE_72_clock = clock;
  assign PE_72_reset = reset;
  assign PE_72_io_data_2_in_bits = PENetwork_32_io_to_pes_9_in_bits; // @[pearray.scala 157:34]
  assign PE_72_io_data_1_in_valid = PENetwork_25_io_to_pes_0_in_valid; // @[pearray.scala 157:34]
  assign PE_72_io_data_1_in_bits = PENetwork_25_io_to_pes_0_in_bits; // @[pearray.scala 157:34]
  assign PE_72_io_data_0_in_valid = 1'h0; // @[pearray.scala 157:34]
  assign PE_72_io_data_0_in_bits = 8'h0; // @[pearray.scala 157:34]
  assign PE_72_io_sig_stat2trans = _T_898_3; // @[pearray.scala 180:38]
  assign PE_73_clock = clock;
  assign PE_73_reset = reset;
  assign PE_73_io_data_2_in_bits = PENetwork_33_io_to_pes_9_in_bits; // @[pearray.scala 157:34]
  assign PE_73_io_data_1_in_valid = PENetwork_25_io_to_pes_1_in_valid; // @[pearray.scala 157:34]
  assign PE_73_io_data_1_in_bits = PENetwork_25_io_to_pes_1_in_bits; // @[pearray.scala 157:34]
  assign PE_73_io_data_0_in_valid = PENetwork_9_io_to_pes_1_in_valid; // @[pearray.scala 157:34]
  assign PE_73_io_data_0_in_bits = PENetwork_9_io_to_pes_1_in_bits; // @[pearray.scala 157:34]
  assign PE_73_io_sig_stat2trans = _T_910_3; // @[pearray.scala 180:38]
  assign PE_74_clock = clock;
  assign PE_74_reset = reset;
  assign PE_74_io_data_2_in_bits = PENetwork_34_io_to_pes_9_in_bits; // @[pearray.scala 157:34]
  assign PE_74_io_data_1_in_valid = PENetwork_25_io_to_pes_2_in_valid; // @[pearray.scala 157:34]
  assign PE_74_io_data_1_in_bits = PENetwork_25_io_to_pes_2_in_bits; // @[pearray.scala 157:34]
  assign PE_74_io_data_0_in_valid = PENetwork_9_io_to_pes_2_in_valid; // @[pearray.scala 157:34]
  assign PE_74_io_data_0_in_bits = PENetwork_9_io_to_pes_2_in_bits; // @[pearray.scala 157:34]
  assign PE_74_io_sig_stat2trans = _T_922_3; // @[pearray.scala 180:38]
  assign PE_75_clock = clock;
  assign PE_75_reset = reset;
  assign PE_75_io_data_2_in_bits = PENetwork_35_io_to_pes_9_in_bits; // @[pearray.scala 157:34]
  assign PE_75_io_data_1_in_valid = PENetwork_25_io_to_pes_3_in_valid; // @[pearray.scala 157:34]
  assign PE_75_io_data_1_in_bits = PENetwork_25_io_to_pes_3_in_bits; // @[pearray.scala 157:34]
  assign PE_75_io_data_0_in_valid = PENetwork_9_io_to_pes_3_in_valid; // @[pearray.scala 157:34]
  assign PE_75_io_data_0_in_bits = PENetwork_9_io_to_pes_3_in_bits; // @[pearray.scala 157:34]
  assign PE_75_io_sig_stat2trans = _T_934_3; // @[pearray.scala 180:38]
  assign PE_76_clock = clock;
  assign PE_76_reset = reset;
  assign PE_76_io_data_2_in_bits = PENetwork_36_io_to_pes_9_in_bits; // @[pearray.scala 157:34]
  assign PE_76_io_data_1_in_valid = PENetwork_25_io_to_pes_4_in_valid; // @[pearray.scala 157:34]
  assign PE_76_io_data_1_in_bits = PENetwork_25_io_to_pes_4_in_bits; // @[pearray.scala 157:34]
  assign PE_76_io_data_0_in_valid = PENetwork_9_io_to_pes_4_in_valid; // @[pearray.scala 157:34]
  assign PE_76_io_data_0_in_bits = PENetwork_9_io_to_pes_4_in_bits; // @[pearray.scala 157:34]
  assign PE_76_io_sig_stat2trans = _T_946_3; // @[pearray.scala 180:38]
  assign PE_77_clock = clock;
  assign PE_77_reset = reset;
  assign PE_77_io_data_2_in_bits = PENetwork_37_io_to_pes_9_in_bits; // @[pearray.scala 157:34]
  assign PE_77_io_data_1_in_valid = PENetwork_25_io_to_pes_5_in_valid; // @[pearray.scala 157:34]
  assign PE_77_io_data_1_in_bits = PENetwork_25_io_to_pes_5_in_bits; // @[pearray.scala 157:34]
  assign PE_77_io_data_0_in_valid = PENetwork_9_io_to_pes_5_in_valid; // @[pearray.scala 157:34]
  assign PE_77_io_data_0_in_bits = PENetwork_9_io_to_pes_5_in_bits; // @[pearray.scala 157:34]
  assign PE_77_io_sig_stat2trans = _T_958_3; // @[pearray.scala 180:38]
  assign PE_78_clock = clock;
  assign PE_78_reset = reset;
  assign PE_78_io_data_2_in_bits = PENetwork_38_io_to_pes_9_in_bits; // @[pearray.scala 157:34]
  assign PE_78_io_data_1_in_valid = PENetwork_25_io_to_pes_6_in_valid; // @[pearray.scala 157:34]
  assign PE_78_io_data_1_in_bits = PENetwork_25_io_to_pes_6_in_bits; // @[pearray.scala 157:34]
  assign PE_78_io_data_0_in_valid = PENetwork_9_io_to_pes_6_in_valid; // @[pearray.scala 157:34]
  assign PE_78_io_data_0_in_bits = PENetwork_9_io_to_pes_6_in_bits; // @[pearray.scala 157:34]
  assign PE_78_io_sig_stat2trans = _T_970_3; // @[pearray.scala 180:38]
  assign PE_79_clock = clock;
  assign PE_79_reset = reset;
  assign PE_79_io_data_2_in_bits = PENetwork_39_io_to_pes_9_in_bits; // @[pearray.scala 157:34]
  assign PE_79_io_data_1_in_valid = PENetwork_25_io_to_pes_7_in_valid; // @[pearray.scala 157:34]
  assign PE_79_io_data_1_in_bits = PENetwork_25_io_to_pes_7_in_bits; // @[pearray.scala 157:34]
  assign PE_79_io_data_0_in_valid = PENetwork_9_io_to_pes_7_in_valid; // @[pearray.scala 157:34]
  assign PE_79_io_data_0_in_bits = PENetwork_9_io_to_pes_7_in_bits; // @[pearray.scala 157:34]
  assign PE_79_io_sig_stat2trans = _T_982_3; // @[pearray.scala 180:38]
  assign PE_80_clock = clock;
  assign PE_80_reset = reset;
  assign PE_80_io_data_2_in_bits = PENetwork_32_io_to_pes_10_in_bits; // @[pearray.scala 157:34]
  assign PE_80_io_data_1_in_valid = PENetwork_26_io_to_pes_0_in_valid; // @[pearray.scala 157:34]
  assign PE_80_io_data_1_in_bits = PENetwork_26_io_to_pes_0_in_bits; // @[pearray.scala 157:34]
  assign PE_80_io_data_0_in_valid = 1'h0; // @[pearray.scala 157:34]
  assign PE_80_io_data_0_in_bits = 8'h0; // @[pearray.scala 157:34]
  assign PE_80_io_sig_stat2trans = _T_996_3; // @[pearray.scala 180:38]
  assign PE_81_clock = clock;
  assign PE_81_reset = reset;
  assign PE_81_io_data_2_in_bits = PENetwork_33_io_to_pes_10_in_bits; // @[pearray.scala 157:34]
  assign PE_81_io_data_1_in_valid = PENetwork_26_io_to_pes_1_in_valid; // @[pearray.scala 157:34]
  assign PE_81_io_data_1_in_bits = PENetwork_26_io_to_pes_1_in_bits; // @[pearray.scala 157:34]
  assign PE_81_io_data_0_in_valid = PENetwork_10_io_to_pes_1_in_valid; // @[pearray.scala 157:34]
  assign PE_81_io_data_0_in_bits = PENetwork_10_io_to_pes_1_in_bits; // @[pearray.scala 157:34]
  assign PE_81_io_sig_stat2trans = _T_1008_3; // @[pearray.scala 180:38]
  assign PE_82_clock = clock;
  assign PE_82_reset = reset;
  assign PE_82_io_data_2_in_bits = PENetwork_34_io_to_pes_10_in_bits; // @[pearray.scala 157:34]
  assign PE_82_io_data_1_in_valid = PENetwork_26_io_to_pes_2_in_valid; // @[pearray.scala 157:34]
  assign PE_82_io_data_1_in_bits = PENetwork_26_io_to_pes_2_in_bits; // @[pearray.scala 157:34]
  assign PE_82_io_data_0_in_valid = PENetwork_10_io_to_pes_2_in_valid; // @[pearray.scala 157:34]
  assign PE_82_io_data_0_in_bits = PENetwork_10_io_to_pes_2_in_bits; // @[pearray.scala 157:34]
  assign PE_82_io_sig_stat2trans = _T_1020_3; // @[pearray.scala 180:38]
  assign PE_83_clock = clock;
  assign PE_83_reset = reset;
  assign PE_83_io_data_2_in_bits = PENetwork_35_io_to_pes_10_in_bits; // @[pearray.scala 157:34]
  assign PE_83_io_data_1_in_valid = PENetwork_26_io_to_pes_3_in_valid; // @[pearray.scala 157:34]
  assign PE_83_io_data_1_in_bits = PENetwork_26_io_to_pes_3_in_bits; // @[pearray.scala 157:34]
  assign PE_83_io_data_0_in_valid = PENetwork_10_io_to_pes_3_in_valid; // @[pearray.scala 157:34]
  assign PE_83_io_data_0_in_bits = PENetwork_10_io_to_pes_3_in_bits; // @[pearray.scala 157:34]
  assign PE_83_io_sig_stat2trans = _T_1032_3; // @[pearray.scala 180:38]
  assign PE_84_clock = clock;
  assign PE_84_reset = reset;
  assign PE_84_io_data_2_in_bits = PENetwork_36_io_to_pes_10_in_bits; // @[pearray.scala 157:34]
  assign PE_84_io_data_1_in_valid = PENetwork_26_io_to_pes_4_in_valid; // @[pearray.scala 157:34]
  assign PE_84_io_data_1_in_bits = PENetwork_26_io_to_pes_4_in_bits; // @[pearray.scala 157:34]
  assign PE_84_io_data_0_in_valid = PENetwork_10_io_to_pes_4_in_valid; // @[pearray.scala 157:34]
  assign PE_84_io_data_0_in_bits = PENetwork_10_io_to_pes_4_in_bits; // @[pearray.scala 157:34]
  assign PE_84_io_sig_stat2trans = _T_1044_3; // @[pearray.scala 180:38]
  assign PE_85_clock = clock;
  assign PE_85_reset = reset;
  assign PE_85_io_data_2_in_bits = PENetwork_37_io_to_pes_10_in_bits; // @[pearray.scala 157:34]
  assign PE_85_io_data_1_in_valid = PENetwork_26_io_to_pes_5_in_valid; // @[pearray.scala 157:34]
  assign PE_85_io_data_1_in_bits = PENetwork_26_io_to_pes_5_in_bits; // @[pearray.scala 157:34]
  assign PE_85_io_data_0_in_valid = PENetwork_10_io_to_pes_5_in_valid; // @[pearray.scala 157:34]
  assign PE_85_io_data_0_in_bits = PENetwork_10_io_to_pes_5_in_bits; // @[pearray.scala 157:34]
  assign PE_85_io_sig_stat2trans = _T_1056_3; // @[pearray.scala 180:38]
  assign PE_86_clock = clock;
  assign PE_86_reset = reset;
  assign PE_86_io_data_2_in_bits = PENetwork_38_io_to_pes_10_in_bits; // @[pearray.scala 157:34]
  assign PE_86_io_data_1_in_valid = PENetwork_26_io_to_pes_6_in_valid; // @[pearray.scala 157:34]
  assign PE_86_io_data_1_in_bits = PENetwork_26_io_to_pes_6_in_bits; // @[pearray.scala 157:34]
  assign PE_86_io_data_0_in_valid = PENetwork_10_io_to_pes_6_in_valid; // @[pearray.scala 157:34]
  assign PE_86_io_data_0_in_bits = PENetwork_10_io_to_pes_6_in_bits; // @[pearray.scala 157:34]
  assign PE_86_io_sig_stat2trans = _T_1068_3; // @[pearray.scala 180:38]
  assign PE_87_clock = clock;
  assign PE_87_reset = reset;
  assign PE_87_io_data_2_in_bits = PENetwork_39_io_to_pes_10_in_bits; // @[pearray.scala 157:34]
  assign PE_87_io_data_1_in_valid = PENetwork_26_io_to_pes_7_in_valid; // @[pearray.scala 157:34]
  assign PE_87_io_data_1_in_bits = PENetwork_26_io_to_pes_7_in_bits; // @[pearray.scala 157:34]
  assign PE_87_io_data_0_in_valid = PENetwork_10_io_to_pes_7_in_valid; // @[pearray.scala 157:34]
  assign PE_87_io_data_0_in_bits = PENetwork_10_io_to_pes_7_in_bits; // @[pearray.scala 157:34]
  assign PE_87_io_sig_stat2trans = _T_1080_3; // @[pearray.scala 180:38]
  assign PE_88_clock = clock;
  assign PE_88_reset = reset;
  assign PE_88_io_data_2_in_bits = PENetwork_32_io_to_pes_11_in_bits; // @[pearray.scala 157:34]
  assign PE_88_io_data_1_in_valid = PENetwork_27_io_to_pes_0_in_valid; // @[pearray.scala 157:34]
  assign PE_88_io_data_1_in_bits = PENetwork_27_io_to_pes_0_in_bits; // @[pearray.scala 157:34]
  assign PE_88_io_data_0_in_valid = 1'h0; // @[pearray.scala 157:34]
  assign PE_88_io_data_0_in_bits = 8'h0; // @[pearray.scala 157:34]
  assign PE_88_io_sig_stat2trans = _T_1094_3; // @[pearray.scala 180:38]
  assign PE_89_clock = clock;
  assign PE_89_reset = reset;
  assign PE_89_io_data_2_in_bits = PENetwork_33_io_to_pes_11_in_bits; // @[pearray.scala 157:34]
  assign PE_89_io_data_1_in_valid = PENetwork_27_io_to_pes_1_in_valid; // @[pearray.scala 157:34]
  assign PE_89_io_data_1_in_bits = PENetwork_27_io_to_pes_1_in_bits; // @[pearray.scala 157:34]
  assign PE_89_io_data_0_in_valid = PENetwork_11_io_to_pes_1_in_valid; // @[pearray.scala 157:34]
  assign PE_89_io_data_0_in_bits = PENetwork_11_io_to_pes_1_in_bits; // @[pearray.scala 157:34]
  assign PE_89_io_sig_stat2trans = _T_1106_3; // @[pearray.scala 180:38]
  assign PE_90_clock = clock;
  assign PE_90_reset = reset;
  assign PE_90_io_data_2_in_bits = PENetwork_34_io_to_pes_11_in_bits; // @[pearray.scala 157:34]
  assign PE_90_io_data_1_in_valid = PENetwork_27_io_to_pes_2_in_valid; // @[pearray.scala 157:34]
  assign PE_90_io_data_1_in_bits = PENetwork_27_io_to_pes_2_in_bits; // @[pearray.scala 157:34]
  assign PE_90_io_data_0_in_valid = PENetwork_11_io_to_pes_2_in_valid; // @[pearray.scala 157:34]
  assign PE_90_io_data_0_in_bits = PENetwork_11_io_to_pes_2_in_bits; // @[pearray.scala 157:34]
  assign PE_90_io_sig_stat2trans = _T_1118_3; // @[pearray.scala 180:38]
  assign PE_91_clock = clock;
  assign PE_91_reset = reset;
  assign PE_91_io_data_2_in_bits = PENetwork_35_io_to_pes_11_in_bits; // @[pearray.scala 157:34]
  assign PE_91_io_data_1_in_valid = PENetwork_27_io_to_pes_3_in_valid; // @[pearray.scala 157:34]
  assign PE_91_io_data_1_in_bits = PENetwork_27_io_to_pes_3_in_bits; // @[pearray.scala 157:34]
  assign PE_91_io_data_0_in_valid = PENetwork_11_io_to_pes_3_in_valid; // @[pearray.scala 157:34]
  assign PE_91_io_data_0_in_bits = PENetwork_11_io_to_pes_3_in_bits; // @[pearray.scala 157:34]
  assign PE_91_io_sig_stat2trans = _T_1130_3; // @[pearray.scala 180:38]
  assign PE_92_clock = clock;
  assign PE_92_reset = reset;
  assign PE_92_io_data_2_in_bits = PENetwork_36_io_to_pes_11_in_bits; // @[pearray.scala 157:34]
  assign PE_92_io_data_1_in_valid = PENetwork_27_io_to_pes_4_in_valid; // @[pearray.scala 157:34]
  assign PE_92_io_data_1_in_bits = PENetwork_27_io_to_pes_4_in_bits; // @[pearray.scala 157:34]
  assign PE_92_io_data_0_in_valid = PENetwork_11_io_to_pes_4_in_valid; // @[pearray.scala 157:34]
  assign PE_92_io_data_0_in_bits = PENetwork_11_io_to_pes_4_in_bits; // @[pearray.scala 157:34]
  assign PE_92_io_sig_stat2trans = _T_1142_3; // @[pearray.scala 180:38]
  assign PE_93_clock = clock;
  assign PE_93_reset = reset;
  assign PE_93_io_data_2_in_bits = PENetwork_37_io_to_pes_11_in_bits; // @[pearray.scala 157:34]
  assign PE_93_io_data_1_in_valid = PENetwork_27_io_to_pes_5_in_valid; // @[pearray.scala 157:34]
  assign PE_93_io_data_1_in_bits = PENetwork_27_io_to_pes_5_in_bits; // @[pearray.scala 157:34]
  assign PE_93_io_data_0_in_valid = PENetwork_11_io_to_pes_5_in_valid; // @[pearray.scala 157:34]
  assign PE_93_io_data_0_in_bits = PENetwork_11_io_to_pes_5_in_bits; // @[pearray.scala 157:34]
  assign PE_93_io_sig_stat2trans = _T_1154_3; // @[pearray.scala 180:38]
  assign PE_94_clock = clock;
  assign PE_94_reset = reset;
  assign PE_94_io_data_2_in_bits = PENetwork_38_io_to_pes_11_in_bits; // @[pearray.scala 157:34]
  assign PE_94_io_data_1_in_valid = PENetwork_27_io_to_pes_6_in_valid; // @[pearray.scala 157:34]
  assign PE_94_io_data_1_in_bits = PENetwork_27_io_to_pes_6_in_bits; // @[pearray.scala 157:34]
  assign PE_94_io_data_0_in_valid = PENetwork_11_io_to_pes_6_in_valid; // @[pearray.scala 157:34]
  assign PE_94_io_data_0_in_bits = PENetwork_11_io_to_pes_6_in_bits; // @[pearray.scala 157:34]
  assign PE_94_io_sig_stat2trans = _T_1166_3; // @[pearray.scala 180:38]
  assign PE_95_clock = clock;
  assign PE_95_reset = reset;
  assign PE_95_io_data_2_in_bits = PENetwork_39_io_to_pes_11_in_bits; // @[pearray.scala 157:34]
  assign PE_95_io_data_1_in_valid = PENetwork_27_io_to_pes_7_in_valid; // @[pearray.scala 157:34]
  assign PE_95_io_data_1_in_bits = PENetwork_27_io_to_pes_7_in_bits; // @[pearray.scala 157:34]
  assign PE_95_io_data_0_in_valid = PENetwork_11_io_to_pes_7_in_valid; // @[pearray.scala 157:34]
  assign PE_95_io_data_0_in_bits = PENetwork_11_io_to_pes_7_in_bits; // @[pearray.scala 157:34]
  assign PE_95_io_sig_stat2trans = _T_1178_3; // @[pearray.scala 180:38]
  assign PE_96_clock = clock;
  assign PE_96_reset = reset;
  assign PE_96_io_data_2_in_bits = PENetwork_32_io_to_pes_12_in_bits; // @[pearray.scala 157:34]
  assign PE_96_io_data_1_in_valid = PENetwork_28_io_to_pes_0_in_valid; // @[pearray.scala 157:34]
  assign PE_96_io_data_1_in_bits = PENetwork_28_io_to_pes_0_in_bits; // @[pearray.scala 157:34]
  assign PE_96_io_data_0_in_valid = 1'h0; // @[pearray.scala 157:34]
  assign PE_96_io_data_0_in_bits = 8'h0; // @[pearray.scala 157:34]
  assign PE_96_io_sig_stat2trans = _T_1192_3; // @[pearray.scala 180:38]
  assign PE_97_clock = clock;
  assign PE_97_reset = reset;
  assign PE_97_io_data_2_in_bits = PENetwork_33_io_to_pes_12_in_bits; // @[pearray.scala 157:34]
  assign PE_97_io_data_1_in_valid = PENetwork_28_io_to_pes_1_in_valid; // @[pearray.scala 157:34]
  assign PE_97_io_data_1_in_bits = PENetwork_28_io_to_pes_1_in_bits; // @[pearray.scala 157:34]
  assign PE_97_io_data_0_in_valid = PENetwork_12_io_to_pes_1_in_valid; // @[pearray.scala 157:34]
  assign PE_97_io_data_0_in_bits = PENetwork_12_io_to_pes_1_in_bits; // @[pearray.scala 157:34]
  assign PE_97_io_sig_stat2trans = _T_1204_3; // @[pearray.scala 180:38]
  assign PE_98_clock = clock;
  assign PE_98_reset = reset;
  assign PE_98_io_data_2_in_bits = PENetwork_34_io_to_pes_12_in_bits; // @[pearray.scala 157:34]
  assign PE_98_io_data_1_in_valid = PENetwork_28_io_to_pes_2_in_valid; // @[pearray.scala 157:34]
  assign PE_98_io_data_1_in_bits = PENetwork_28_io_to_pes_2_in_bits; // @[pearray.scala 157:34]
  assign PE_98_io_data_0_in_valid = PENetwork_12_io_to_pes_2_in_valid; // @[pearray.scala 157:34]
  assign PE_98_io_data_0_in_bits = PENetwork_12_io_to_pes_2_in_bits; // @[pearray.scala 157:34]
  assign PE_98_io_sig_stat2trans = _T_1216_3; // @[pearray.scala 180:38]
  assign PE_99_clock = clock;
  assign PE_99_reset = reset;
  assign PE_99_io_data_2_in_bits = PENetwork_35_io_to_pes_12_in_bits; // @[pearray.scala 157:34]
  assign PE_99_io_data_1_in_valid = PENetwork_28_io_to_pes_3_in_valid; // @[pearray.scala 157:34]
  assign PE_99_io_data_1_in_bits = PENetwork_28_io_to_pes_3_in_bits; // @[pearray.scala 157:34]
  assign PE_99_io_data_0_in_valid = PENetwork_12_io_to_pes_3_in_valid; // @[pearray.scala 157:34]
  assign PE_99_io_data_0_in_bits = PENetwork_12_io_to_pes_3_in_bits; // @[pearray.scala 157:34]
  assign PE_99_io_sig_stat2trans = _T_1228_3; // @[pearray.scala 180:38]
  assign PE_100_clock = clock;
  assign PE_100_reset = reset;
  assign PE_100_io_data_2_in_bits = PENetwork_36_io_to_pes_12_in_bits; // @[pearray.scala 157:34]
  assign PE_100_io_data_1_in_valid = PENetwork_28_io_to_pes_4_in_valid; // @[pearray.scala 157:34]
  assign PE_100_io_data_1_in_bits = PENetwork_28_io_to_pes_4_in_bits; // @[pearray.scala 157:34]
  assign PE_100_io_data_0_in_valid = PENetwork_12_io_to_pes_4_in_valid; // @[pearray.scala 157:34]
  assign PE_100_io_data_0_in_bits = PENetwork_12_io_to_pes_4_in_bits; // @[pearray.scala 157:34]
  assign PE_100_io_sig_stat2trans = _T_1240_3; // @[pearray.scala 180:38]
  assign PE_101_clock = clock;
  assign PE_101_reset = reset;
  assign PE_101_io_data_2_in_bits = PENetwork_37_io_to_pes_12_in_bits; // @[pearray.scala 157:34]
  assign PE_101_io_data_1_in_valid = PENetwork_28_io_to_pes_5_in_valid; // @[pearray.scala 157:34]
  assign PE_101_io_data_1_in_bits = PENetwork_28_io_to_pes_5_in_bits; // @[pearray.scala 157:34]
  assign PE_101_io_data_0_in_valid = PENetwork_12_io_to_pes_5_in_valid; // @[pearray.scala 157:34]
  assign PE_101_io_data_0_in_bits = PENetwork_12_io_to_pes_5_in_bits; // @[pearray.scala 157:34]
  assign PE_101_io_sig_stat2trans = _T_1252_3; // @[pearray.scala 180:38]
  assign PE_102_clock = clock;
  assign PE_102_reset = reset;
  assign PE_102_io_data_2_in_bits = PENetwork_38_io_to_pes_12_in_bits; // @[pearray.scala 157:34]
  assign PE_102_io_data_1_in_valid = PENetwork_28_io_to_pes_6_in_valid; // @[pearray.scala 157:34]
  assign PE_102_io_data_1_in_bits = PENetwork_28_io_to_pes_6_in_bits; // @[pearray.scala 157:34]
  assign PE_102_io_data_0_in_valid = PENetwork_12_io_to_pes_6_in_valid; // @[pearray.scala 157:34]
  assign PE_102_io_data_0_in_bits = PENetwork_12_io_to_pes_6_in_bits; // @[pearray.scala 157:34]
  assign PE_102_io_sig_stat2trans = _T_1264_3; // @[pearray.scala 180:38]
  assign PE_103_clock = clock;
  assign PE_103_reset = reset;
  assign PE_103_io_data_2_in_bits = PENetwork_39_io_to_pes_12_in_bits; // @[pearray.scala 157:34]
  assign PE_103_io_data_1_in_valid = PENetwork_28_io_to_pes_7_in_valid; // @[pearray.scala 157:34]
  assign PE_103_io_data_1_in_bits = PENetwork_28_io_to_pes_7_in_bits; // @[pearray.scala 157:34]
  assign PE_103_io_data_0_in_valid = PENetwork_12_io_to_pes_7_in_valid; // @[pearray.scala 157:34]
  assign PE_103_io_data_0_in_bits = PENetwork_12_io_to_pes_7_in_bits; // @[pearray.scala 157:34]
  assign PE_103_io_sig_stat2trans = _T_1276_3; // @[pearray.scala 180:38]
  assign PE_104_clock = clock;
  assign PE_104_reset = reset;
  assign PE_104_io_data_2_in_bits = PENetwork_32_io_to_pes_13_in_bits; // @[pearray.scala 157:34]
  assign PE_104_io_data_1_in_valid = PENetwork_29_io_to_pes_0_in_valid; // @[pearray.scala 157:34]
  assign PE_104_io_data_1_in_bits = PENetwork_29_io_to_pes_0_in_bits; // @[pearray.scala 157:34]
  assign PE_104_io_data_0_in_valid = 1'h0; // @[pearray.scala 157:34]
  assign PE_104_io_data_0_in_bits = 8'h0; // @[pearray.scala 157:34]
  assign PE_104_io_sig_stat2trans = _T_1290_3; // @[pearray.scala 180:38]
  assign PE_105_clock = clock;
  assign PE_105_reset = reset;
  assign PE_105_io_data_2_in_bits = PENetwork_33_io_to_pes_13_in_bits; // @[pearray.scala 157:34]
  assign PE_105_io_data_1_in_valid = PENetwork_29_io_to_pes_1_in_valid; // @[pearray.scala 157:34]
  assign PE_105_io_data_1_in_bits = PENetwork_29_io_to_pes_1_in_bits; // @[pearray.scala 157:34]
  assign PE_105_io_data_0_in_valid = PENetwork_13_io_to_pes_1_in_valid; // @[pearray.scala 157:34]
  assign PE_105_io_data_0_in_bits = PENetwork_13_io_to_pes_1_in_bits; // @[pearray.scala 157:34]
  assign PE_105_io_sig_stat2trans = _T_1302_3; // @[pearray.scala 180:38]
  assign PE_106_clock = clock;
  assign PE_106_reset = reset;
  assign PE_106_io_data_2_in_bits = PENetwork_34_io_to_pes_13_in_bits; // @[pearray.scala 157:34]
  assign PE_106_io_data_1_in_valid = PENetwork_29_io_to_pes_2_in_valid; // @[pearray.scala 157:34]
  assign PE_106_io_data_1_in_bits = PENetwork_29_io_to_pes_2_in_bits; // @[pearray.scala 157:34]
  assign PE_106_io_data_0_in_valid = PENetwork_13_io_to_pes_2_in_valid; // @[pearray.scala 157:34]
  assign PE_106_io_data_0_in_bits = PENetwork_13_io_to_pes_2_in_bits; // @[pearray.scala 157:34]
  assign PE_106_io_sig_stat2trans = _T_1314_3; // @[pearray.scala 180:38]
  assign PE_107_clock = clock;
  assign PE_107_reset = reset;
  assign PE_107_io_data_2_in_bits = PENetwork_35_io_to_pes_13_in_bits; // @[pearray.scala 157:34]
  assign PE_107_io_data_1_in_valid = PENetwork_29_io_to_pes_3_in_valid; // @[pearray.scala 157:34]
  assign PE_107_io_data_1_in_bits = PENetwork_29_io_to_pes_3_in_bits; // @[pearray.scala 157:34]
  assign PE_107_io_data_0_in_valid = PENetwork_13_io_to_pes_3_in_valid; // @[pearray.scala 157:34]
  assign PE_107_io_data_0_in_bits = PENetwork_13_io_to_pes_3_in_bits; // @[pearray.scala 157:34]
  assign PE_107_io_sig_stat2trans = _T_1326_3; // @[pearray.scala 180:38]
  assign PE_108_clock = clock;
  assign PE_108_reset = reset;
  assign PE_108_io_data_2_in_bits = PENetwork_36_io_to_pes_13_in_bits; // @[pearray.scala 157:34]
  assign PE_108_io_data_1_in_valid = PENetwork_29_io_to_pes_4_in_valid; // @[pearray.scala 157:34]
  assign PE_108_io_data_1_in_bits = PENetwork_29_io_to_pes_4_in_bits; // @[pearray.scala 157:34]
  assign PE_108_io_data_0_in_valid = PENetwork_13_io_to_pes_4_in_valid; // @[pearray.scala 157:34]
  assign PE_108_io_data_0_in_bits = PENetwork_13_io_to_pes_4_in_bits; // @[pearray.scala 157:34]
  assign PE_108_io_sig_stat2trans = _T_1338_3; // @[pearray.scala 180:38]
  assign PE_109_clock = clock;
  assign PE_109_reset = reset;
  assign PE_109_io_data_2_in_bits = PENetwork_37_io_to_pes_13_in_bits; // @[pearray.scala 157:34]
  assign PE_109_io_data_1_in_valid = PENetwork_29_io_to_pes_5_in_valid; // @[pearray.scala 157:34]
  assign PE_109_io_data_1_in_bits = PENetwork_29_io_to_pes_5_in_bits; // @[pearray.scala 157:34]
  assign PE_109_io_data_0_in_valid = PENetwork_13_io_to_pes_5_in_valid; // @[pearray.scala 157:34]
  assign PE_109_io_data_0_in_bits = PENetwork_13_io_to_pes_5_in_bits; // @[pearray.scala 157:34]
  assign PE_109_io_sig_stat2trans = _T_1350_3; // @[pearray.scala 180:38]
  assign PE_110_clock = clock;
  assign PE_110_reset = reset;
  assign PE_110_io_data_2_in_bits = PENetwork_38_io_to_pes_13_in_bits; // @[pearray.scala 157:34]
  assign PE_110_io_data_1_in_valid = PENetwork_29_io_to_pes_6_in_valid; // @[pearray.scala 157:34]
  assign PE_110_io_data_1_in_bits = PENetwork_29_io_to_pes_6_in_bits; // @[pearray.scala 157:34]
  assign PE_110_io_data_0_in_valid = PENetwork_13_io_to_pes_6_in_valid; // @[pearray.scala 157:34]
  assign PE_110_io_data_0_in_bits = PENetwork_13_io_to_pes_6_in_bits; // @[pearray.scala 157:34]
  assign PE_110_io_sig_stat2trans = _T_1362_3; // @[pearray.scala 180:38]
  assign PE_111_clock = clock;
  assign PE_111_reset = reset;
  assign PE_111_io_data_2_in_bits = PENetwork_39_io_to_pes_13_in_bits; // @[pearray.scala 157:34]
  assign PE_111_io_data_1_in_valid = PENetwork_29_io_to_pes_7_in_valid; // @[pearray.scala 157:34]
  assign PE_111_io_data_1_in_bits = PENetwork_29_io_to_pes_7_in_bits; // @[pearray.scala 157:34]
  assign PE_111_io_data_0_in_valid = PENetwork_13_io_to_pes_7_in_valid; // @[pearray.scala 157:34]
  assign PE_111_io_data_0_in_bits = PENetwork_13_io_to_pes_7_in_bits; // @[pearray.scala 157:34]
  assign PE_111_io_sig_stat2trans = _T_1374_3; // @[pearray.scala 180:38]
  assign PE_112_clock = clock;
  assign PE_112_reset = reset;
  assign PE_112_io_data_2_in_bits = PENetwork_32_io_to_pes_14_in_bits; // @[pearray.scala 157:34]
  assign PE_112_io_data_1_in_valid = PENetwork_30_io_to_pes_0_in_valid; // @[pearray.scala 157:34]
  assign PE_112_io_data_1_in_bits = PENetwork_30_io_to_pes_0_in_bits; // @[pearray.scala 157:34]
  assign PE_112_io_data_0_in_valid = 1'h0; // @[pearray.scala 157:34]
  assign PE_112_io_data_0_in_bits = 8'h0; // @[pearray.scala 157:34]
  assign PE_112_io_sig_stat2trans = _T_1388_3; // @[pearray.scala 180:38]
  assign PE_113_clock = clock;
  assign PE_113_reset = reset;
  assign PE_113_io_data_2_in_bits = PENetwork_33_io_to_pes_14_in_bits; // @[pearray.scala 157:34]
  assign PE_113_io_data_1_in_valid = PENetwork_30_io_to_pes_1_in_valid; // @[pearray.scala 157:34]
  assign PE_113_io_data_1_in_bits = PENetwork_30_io_to_pes_1_in_bits; // @[pearray.scala 157:34]
  assign PE_113_io_data_0_in_valid = PENetwork_14_io_to_pes_1_in_valid; // @[pearray.scala 157:34]
  assign PE_113_io_data_0_in_bits = PENetwork_14_io_to_pes_1_in_bits; // @[pearray.scala 157:34]
  assign PE_113_io_sig_stat2trans = _T_1400_3; // @[pearray.scala 180:38]
  assign PE_114_clock = clock;
  assign PE_114_reset = reset;
  assign PE_114_io_data_2_in_bits = PENetwork_34_io_to_pes_14_in_bits; // @[pearray.scala 157:34]
  assign PE_114_io_data_1_in_valid = PENetwork_30_io_to_pes_2_in_valid; // @[pearray.scala 157:34]
  assign PE_114_io_data_1_in_bits = PENetwork_30_io_to_pes_2_in_bits; // @[pearray.scala 157:34]
  assign PE_114_io_data_0_in_valid = PENetwork_14_io_to_pes_2_in_valid; // @[pearray.scala 157:34]
  assign PE_114_io_data_0_in_bits = PENetwork_14_io_to_pes_2_in_bits; // @[pearray.scala 157:34]
  assign PE_114_io_sig_stat2trans = _T_1412_3; // @[pearray.scala 180:38]
  assign PE_115_clock = clock;
  assign PE_115_reset = reset;
  assign PE_115_io_data_2_in_bits = PENetwork_35_io_to_pes_14_in_bits; // @[pearray.scala 157:34]
  assign PE_115_io_data_1_in_valid = PENetwork_30_io_to_pes_3_in_valid; // @[pearray.scala 157:34]
  assign PE_115_io_data_1_in_bits = PENetwork_30_io_to_pes_3_in_bits; // @[pearray.scala 157:34]
  assign PE_115_io_data_0_in_valid = PENetwork_14_io_to_pes_3_in_valid; // @[pearray.scala 157:34]
  assign PE_115_io_data_0_in_bits = PENetwork_14_io_to_pes_3_in_bits; // @[pearray.scala 157:34]
  assign PE_115_io_sig_stat2trans = _T_1424_3; // @[pearray.scala 180:38]
  assign PE_116_clock = clock;
  assign PE_116_reset = reset;
  assign PE_116_io_data_2_in_bits = PENetwork_36_io_to_pes_14_in_bits; // @[pearray.scala 157:34]
  assign PE_116_io_data_1_in_valid = PENetwork_30_io_to_pes_4_in_valid; // @[pearray.scala 157:34]
  assign PE_116_io_data_1_in_bits = PENetwork_30_io_to_pes_4_in_bits; // @[pearray.scala 157:34]
  assign PE_116_io_data_0_in_valid = PENetwork_14_io_to_pes_4_in_valid; // @[pearray.scala 157:34]
  assign PE_116_io_data_0_in_bits = PENetwork_14_io_to_pes_4_in_bits; // @[pearray.scala 157:34]
  assign PE_116_io_sig_stat2trans = _T_1436_3; // @[pearray.scala 180:38]
  assign PE_117_clock = clock;
  assign PE_117_reset = reset;
  assign PE_117_io_data_2_in_bits = PENetwork_37_io_to_pes_14_in_bits; // @[pearray.scala 157:34]
  assign PE_117_io_data_1_in_valid = PENetwork_30_io_to_pes_5_in_valid; // @[pearray.scala 157:34]
  assign PE_117_io_data_1_in_bits = PENetwork_30_io_to_pes_5_in_bits; // @[pearray.scala 157:34]
  assign PE_117_io_data_0_in_valid = PENetwork_14_io_to_pes_5_in_valid; // @[pearray.scala 157:34]
  assign PE_117_io_data_0_in_bits = PENetwork_14_io_to_pes_5_in_bits; // @[pearray.scala 157:34]
  assign PE_117_io_sig_stat2trans = _T_1448_3; // @[pearray.scala 180:38]
  assign PE_118_clock = clock;
  assign PE_118_reset = reset;
  assign PE_118_io_data_2_in_bits = PENetwork_38_io_to_pes_14_in_bits; // @[pearray.scala 157:34]
  assign PE_118_io_data_1_in_valid = PENetwork_30_io_to_pes_6_in_valid; // @[pearray.scala 157:34]
  assign PE_118_io_data_1_in_bits = PENetwork_30_io_to_pes_6_in_bits; // @[pearray.scala 157:34]
  assign PE_118_io_data_0_in_valid = PENetwork_14_io_to_pes_6_in_valid; // @[pearray.scala 157:34]
  assign PE_118_io_data_0_in_bits = PENetwork_14_io_to_pes_6_in_bits; // @[pearray.scala 157:34]
  assign PE_118_io_sig_stat2trans = _T_1460_3; // @[pearray.scala 180:38]
  assign PE_119_clock = clock;
  assign PE_119_reset = reset;
  assign PE_119_io_data_2_in_bits = PENetwork_39_io_to_pes_14_in_bits; // @[pearray.scala 157:34]
  assign PE_119_io_data_1_in_valid = PENetwork_30_io_to_pes_7_in_valid; // @[pearray.scala 157:34]
  assign PE_119_io_data_1_in_bits = PENetwork_30_io_to_pes_7_in_bits; // @[pearray.scala 157:34]
  assign PE_119_io_data_0_in_valid = PENetwork_14_io_to_pes_7_in_valid; // @[pearray.scala 157:34]
  assign PE_119_io_data_0_in_bits = PENetwork_14_io_to_pes_7_in_bits; // @[pearray.scala 157:34]
  assign PE_119_io_sig_stat2trans = _T_1472_3; // @[pearray.scala 180:38]
  assign PE_120_clock = clock;
  assign PE_120_reset = reset;
  assign PE_120_io_data_2_in_bits = PENetwork_32_io_to_pes_15_in_bits; // @[pearray.scala 157:34]
  assign PE_120_io_data_1_in_valid = PENetwork_31_io_to_pes_0_in_valid; // @[pearray.scala 157:34]
  assign PE_120_io_data_1_in_bits = PENetwork_31_io_to_pes_0_in_bits; // @[pearray.scala 157:34]
  assign PE_120_io_data_0_in_valid = 1'h0; // @[pearray.scala 157:34]
  assign PE_120_io_data_0_in_bits = 8'h0; // @[pearray.scala 157:34]
  assign PE_120_io_sig_stat2trans = _T_1486_3; // @[pearray.scala 180:38]
  assign PE_121_clock = clock;
  assign PE_121_reset = reset;
  assign PE_121_io_data_2_in_bits = PENetwork_33_io_to_pes_15_in_bits; // @[pearray.scala 157:34]
  assign PE_121_io_data_1_in_valid = PENetwork_31_io_to_pes_1_in_valid; // @[pearray.scala 157:34]
  assign PE_121_io_data_1_in_bits = PENetwork_31_io_to_pes_1_in_bits; // @[pearray.scala 157:34]
  assign PE_121_io_data_0_in_valid = PENetwork_15_io_to_pes_1_in_valid; // @[pearray.scala 157:34]
  assign PE_121_io_data_0_in_bits = PENetwork_15_io_to_pes_1_in_bits; // @[pearray.scala 157:34]
  assign PE_121_io_sig_stat2trans = _T_1498_3; // @[pearray.scala 180:38]
  assign PE_122_clock = clock;
  assign PE_122_reset = reset;
  assign PE_122_io_data_2_in_bits = PENetwork_34_io_to_pes_15_in_bits; // @[pearray.scala 157:34]
  assign PE_122_io_data_1_in_valid = PENetwork_31_io_to_pes_2_in_valid; // @[pearray.scala 157:34]
  assign PE_122_io_data_1_in_bits = PENetwork_31_io_to_pes_2_in_bits; // @[pearray.scala 157:34]
  assign PE_122_io_data_0_in_valid = PENetwork_15_io_to_pes_2_in_valid; // @[pearray.scala 157:34]
  assign PE_122_io_data_0_in_bits = PENetwork_15_io_to_pes_2_in_bits; // @[pearray.scala 157:34]
  assign PE_122_io_sig_stat2trans = _T_1510_3; // @[pearray.scala 180:38]
  assign PE_123_clock = clock;
  assign PE_123_reset = reset;
  assign PE_123_io_data_2_in_bits = PENetwork_35_io_to_pes_15_in_bits; // @[pearray.scala 157:34]
  assign PE_123_io_data_1_in_valid = PENetwork_31_io_to_pes_3_in_valid; // @[pearray.scala 157:34]
  assign PE_123_io_data_1_in_bits = PENetwork_31_io_to_pes_3_in_bits; // @[pearray.scala 157:34]
  assign PE_123_io_data_0_in_valid = PENetwork_15_io_to_pes_3_in_valid; // @[pearray.scala 157:34]
  assign PE_123_io_data_0_in_bits = PENetwork_15_io_to_pes_3_in_bits; // @[pearray.scala 157:34]
  assign PE_123_io_sig_stat2trans = _T_1522_3; // @[pearray.scala 180:38]
  assign PE_124_clock = clock;
  assign PE_124_reset = reset;
  assign PE_124_io_data_2_in_bits = PENetwork_36_io_to_pes_15_in_bits; // @[pearray.scala 157:34]
  assign PE_124_io_data_1_in_valid = PENetwork_31_io_to_pes_4_in_valid; // @[pearray.scala 157:34]
  assign PE_124_io_data_1_in_bits = PENetwork_31_io_to_pes_4_in_bits; // @[pearray.scala 157:34]
  assign PE_124_io_data_0_in_valid = PENetwork_15_io_to_pes_4_in_valid; // @[pearray.scala 157:34]
  assign PE_124_io_data_0_in_bits = PENetwork_15_io_to_pes_4_in_bits; // @[pearray.scala 157:34]
  assign PE_124_io_sig_stat2trans = _T_1534_3; // @[pearray.scala 180:38]
  assign PE_125_clock = clock;
  assign PE_125_reset = reset;
  assign PE_125_io_data_2_in_bits = PENetwork_37_io_to_pes_15_in_bits; // @[pearray.scala 157:34]
  assign PE_125_io_data_1_in_valid = PENetwork_31_io_to_pes_5_in_valid; // @[pearray.scala 157:34]
  assign PE_125_io_data_1_in_bits = PENetwork_31_io_to_pes_5_in_bits; // @[pearray.scala 157:34]
  assign PE_125_io_data_0_in_valid = PENetwork_15_io_to_pes_5_in_valid; // @[pearray.scala 157:34]
  assign PE_125_io_data_0_in_bits = PENetwork_15_io_to_pes_5_in_bits; // @[pearray.scala 157:34]
  assign PE_125_io_sig_stat2trans = _T_1546_3; // @[pearray.scala 180:38]
  assign PE_126_clock = clock;
  assign PE_126_reset = reset;
  assign PE_126_io_data_2_in_bits = PENetwork_38_io_to_pes_15_in_bits; // @[pearray.scala 157:34]
  assign PE_126_io_data_1_in_valid = PENetwork_31_io_to_pes_6_in_valid; // @[pearray.scala 157:34]
  assign PE_126_io_data_1_in_bits = PENetwork_31_io_to_pes_6_in_bits; // @[pearray.scala 157:34]
  assign PE_126_io_data_0_in_valid = PENetwork_15_io_to_pes_6_in_valid; // @[pearray.scala 157:34]
  assign PE_126_io_data_0_in_bits = PENetwork_15_io_to_pes_6_in_bits; // @[pearray.scala 157:34]
  assign PE_126_io_sig_stat2trans = _T_1558_3; // @[pearray.scala 180:38]
  assign PE_127_clock = clock;
  assign PE_127_reset = reset;
  assign PE_127_io_data_2_in_bits = PENetwork_39_io_to_pes_15_in_bits; // @[pearray.scala 157:34]
  assign PE_127_io_data_1_in_valid = PENetwork_31_io_to_pes_7_in_valid; // @[pearray.scala 157:34]
  assign PE_127_io_data_1_in_bits = PENetwork_31_io_to_pes_7_in_bits; // @[pearray.scala 157:34]
  assign PE_127_io_data_0_in_valid = PENetwork_15_io_to_pes_7_in_valid; // @[pearray.scala 157:34]
  assign PE_127_io_data_0_in_bits = PENetwork_15_io_to_pes_7_in_bits; // @[pearray.scala 157:34]
  assign PE_127_io_sig_stat2trans = _T_1570_3; // @[pearray.scala 180:38]
  assign PENetwork_io_to_pes_0_out_valid = PE_io_data_0_out_valid; // @[pearray.scala 156:36]
  assign PENetwork_io_to_pes_0_out_bits = PE_io_data_0_out_bits; // @[pearray.scala 156:36]
  assign PENetwork_io_to_pes_1_out_valid = PE_1_io_data_0_out_valid; // @[pearray.scala 156:36]
  assign PENetwork_io_to_pes_1_out_bits = PE_1_io_data_0_out_bits; // @[pearray.scala 156:36]
  assign PENetwork_io_to_pes_2_out_valid = PE_2_io_data_0_out_valid; // @[pearray.scala 156:36]
  assign PENetwork_io_to_pes_2_out_bits = PE_2_io_data_0_out_bits; // @[pearray.scala 156:36]
  assign PENetwork_io_to_pes_3_out_valid = PE_3_io_data_0_out_valid; // @[pearray.scala 156:36]
  assign PENetwork_io_to_pes_3_out_bits = PE_3_io_data_0_out_bits; // @[pearray.scala 156:36]
  assign PENetwork_io_to_pes_4_out_valid = PE_4_io_data_0_out_valid; // @[pearray.scala 156:36]
  assign PENetwork_io_to_pes_4_out_bits = PE_4_io_data_0_out_bits; // @[pearray.scala 156:36]
  assign PENetwork_io_to_pes_5_out_valid = PE_5_io_data_0_out_valid; // @[pearray.scala 156:36]
  assign PENetwork_io_to_pes_5_out_bits = PE_5_io_data_0_out_bits; // @[pearray.scala 156:36]
  assign PENetwork_io_to_pes_6_out_valid = PE_6_io_data_0_out_valid; // @[pearray.scala 156:36]
  assign PENetwork_io_to_pes_6_out_bits = PE_6_io_data_0_out_bits; // @[pearray.scala 156:36]
  assign PENetwork_io_to_pes_7_out_valid = PE_7_io_data_0_out_valid; // @[pearray.scala 156:36]
  assign PENetwork_io_to_pes_7_out_bits = PE_7_io_data_0_out_bits; // @[pearray.scala 156:36]
  assign PENetwork_1_io_to_pes_0_out_valid = PE_8_io_data_0_out_valid; // @[pearray.scala 156:36]
  assign PENetwork_1_io_to_pes_0_out_bits = PE_8_io_data_0_out_bits; // @[pearray.scala 156:36]
  assign PENetwork_1_io_to_pes_1_out_valid = PE_9_io_data_0_out_valid; // @[pearray.scala 156:36]
  assign PENetwork_1_io_to_pes_1_out_bits = PE_9_io_data_0_out_bits; // @[pearray.scala 156:36]
  assign PENetwork_1_io_to_pes_2_out_valid = PE_10_io_data_0_out_valid; // @[pearray.scala 156:36]
  assign PENetwork_1_io_to_pes_2_out_bits = PE_10_io_data_0_out_bits; // @[pearray.scala 156:36]
  assign PENetwork_1_io_to_pes_3_out_valid = PE_11_io_data_0_out_valid; // @[pearray.scala 156:36]
  assign PENetwork_1_io_to_pes_3_out_bits = PE_11_io_data_0_out_bits; // @[pearray.scala 156:36]
  assign PENetwork_1_io_to_pes_4_out_valid = PE_12_io_data_0_out_valid; // @[pearray.scala 156:36]
  assign PENetwork_1_io_to_pes_4_out_bits = PE_12_io_data_0_out_bits; // @[pearray.scala 156:36]
  assign PENetwork_1_io_to_pes_5_out_valid = PE_13_io_data_0_out_valid; // @[pearray.scala 156:36]
  assign PENetwork_1_io_to_pes_5_out_bits = PE_13_io_data_0_out_bits; // @[pearray.scala 156:36]
  assign PENetwork_1_io_to_pes_6_out_valid = PE_14_io_data_0_out_valid; // @[pearray.scala 156:36]
  assign PENetwork_1_io_to_pes_6_out_bits = PE_14_io_data_0_out_bits; // @[pearray.scala 156:36]
  assign PENetwork_1_io_to_pes_7_out_valid = PE_15_io_data_0_out_valid; // @[pearray.scala 156:36]
  assign PENetwork_1_io_to_pes_7_out_bits = PE_15_io_data_0_out_bits; // @[pearray.scala 156:36]
  assign PENetwork_2_io_to_pes_0_out_valid = PE_16_io_data_0_out_valid; // @[pearray.scala 156:36]
  assign PENetwork_2_io_to_pes_0_out_bits = PE_16_io_data_0_out_bits; // @[pearray.scala 156:36]
  assign PENetwork_2_io_to_pes_1_out_valid = PE_17_io_data_0_out_valid; // @[pearray.scala 156:36]
  assign PENetwork_2_io_to_pes_1_out_bits = PE_17_io_data_0_out_bits; // @[pearray.scala 156:36]
  assign PENetwork_2_io_to_pes_2_out_valid = PE_18_io_data_0_out_valid; // @[pearray.scala 156:36]
  assign PENetwork_2_io_to_pes_2_out_bits = PE_18_io_data_0_out_bits; // @[pearray.scala 156:36]
  assign PENetwork_2_io_to_pes_3_out_valid = PE_19_io_data_0_out_valid; // @[pearray.scala 156:36]
  assign PENetwork_2_io_to_pes_3_out_bits = PE_19_io_data_0_out_bits; // @[pearray.scala 156:36]
  assign PENetwork_2_io_to_pes_4_out_valid = PE_20_io_data_0_out_valid; // @[pearray.scala 156:36]
  assign PENetwork_2_io_to_pes_4_out_bits = PE_20_io_data_0_out_bits; // @[pearray.scala 156:36]
  assign PENetwork_2_io_to_pes_5_out_valid = PE_21_io_data_0_out_valid; // @[pearray.scala 156:36]
  assign PENetwork_2_io_to_pes_5_out_bits = PE_21_io_data_0_out_bits; // @[pearray.scala 156:36]
  assign PENetwork_2_io_to_pes_6_out_valid = PE_22_io_data_0_out_valid; // @[pearray.scala 156:36]
  assign PENetwork_2_io_to_pes_6_out_bits = PE_22_io_data_0_out_bits; // @[pearray.scala 156:36]
  assign PENetwork_2_io_to_pes_7_out_valid = PE_23_io_data_0_out_valid; // @[pearray.scala 156:36]
  assign PENetwork_2_io_to_pes_7_out_bits = PE_23_io_data_0_out_bits; // @[pearray.scala 156:36]
  assign PENetwork_3_io_to_pes_0_out_valid = PE_24_io_data_0_out_valid; // @[pearray.scala 156:36]
  assign PENetwork_3_io_to_pes_0_out_bits = PE_24_io_data_0_out_bits; // @[pearray.scala 156:36]
  assign PENetwork_3_io_to_pes_1_out_valid = PE_25_io_data_0_out_valid; // @[pearray.scala 156:36]
  assign PENetwork_3_io_to_pes_1_out_bits = PE_25_io_data_0_out_bits; // @[pearray.scala 156:36]
  assign PENetwork_3_io_to_pes_2_out_valid = PE_26_io_data_0_out_valid; // @[pearray.scala 156:36]
  assign PENetwork_3_io_to_pes_2_out_bits = PE_26_io_data_0_out_bits; // @[pearray.scala 156:36]
  assign PENetwork_3_io_to_pes_3_out_valid = PE_27_io_data_0_out_valid; // @[pearray.scala 156:36]
  assign PENetwork_3_io_to_pes_3_out_bits = PE_27_io_data_0_out_bits; // @[pearray.scala 156:36]
  assign PENetwork_3_io_to_pes_4_out_valid = PE_28_io_data_0_out_valid; // @[pearray.scala 156:36]
  assign PENetwork_3_io_to_pes_4_out_bits = PE_28_io_data_0_out_bits; // @[pearray.scala 156:36]
  assign PENetwork_3_io_to_pes_5_out_valid = PE_29_io_data_0_out_valid; // @[pearray.scala 156:36]
  assign PENetwork_3_io_to_pes_5_out_bits = PE_29_io_data_0_out_bits; // @[pearray.scala 156:36]
  assign PENetwork_3_io_to_pes_6_out_valid = PE_30_io_data_0_out_valid; // @[pearray.scala 156:36]
  assign PENetwork_3_io_to_pes_6_out_bits = PE_30_io_data_0_out_bits; // @[pearray.scala 156:36]
  assign PENetwork_3_io_to_pes_7_out_valid = PE_31_io_data_0_out_valid; // @[pearray.scala 156:36]
  assign PENetwork_3_io_to_pes_7_out_bits = PE_31_io_data_0_out_bits; // @[pearray.scala 156:36]
  assign PENetwork_4_io_to_pes_0_out_valid = PE_32_io_data_0_out_valid; // @[pearray.scala 156:36]
  assign PENetwork_4_io_to_pes_0_out_bits = PE_32_io_data_0_out_bits; // @[pearray.scala 156:36]
  assign PENetwork_4_io_to_pes_1_out_valid = PE_33_io_data_0_out_valid; // @[pearray.scala 156:36]
  assign PENetwork_4_io_to_pes_1_out_bits = PE_33_io_data_0_out_bits; // @[pearray.scala 156:36]
  assign PENetwork_4_io_to_pes_2_out_valid = PE_34_io_data_0_out_valid; // @[pearray.scala 156:36]
  assign PENetwork_4_io_to_pes_2_out_bits = PE_34_io_data_0_out_bits; // @[pearray.scala 156:36]
  assign PENetwork_4_io_to_pes_3_out_valid = PE_35_io_data_0_out_valid; // @[pearray.scala 156:36]
  assign PENetwork_4_io_to_pes_3_out_bits = PE_35_io_data_0_out_bits; // @[pearray.scala 156:36]
  assign PENetwork_4_io_to_pes_4_out_valid = PE_36_io_data_0_out_valid; // @[pearray.scala 156:36]
  assign PENetwork_4_io_to_pes_4_out_bits = PE_36_io_data_0_out_bits; // @[pearray.scala 156:36]
  assign PENetwork_4_io_to_pes_5_out_valid = PE_37_io_data_0_out_valid; // @[pearray.scala 156:36]
  assign PENetwork_4_io_to_pes_5_out_bits = PE_37_io_data_0_out_bits; // @[pearray.scala 156:36]
  assign PENetwork_4_io_to_pes_6_out_valid = PE_38_io_data_0_out_valid; // @[pearray.scala 156:36]
  assign PENetwork_4_io_to_pes_6_out_bits = PE_38_io_data_0_out_bits; // @[pearray.scala 156:36]
  assign PENetwork_4_io_to_pes_7_out_valid = PE_39_io_data_0_out_valid; // @[pearray.scala 156:36]
  assign PENetwork_4_io_to_pes_7_out_bits = PE_39_io_data_0_out_bits; // @[pearray.scala 156:36]
  assign PENetwork_5_io_to_pes_0_out_valid = PE_40_io_data_0_out_valid; // @[pearray.scala 156:36]
  assign PENetwork_5_io_to_pes_0_out_bits = PE_40_io_data_0_out_bits; // @[pearray.scala 156:36]
  assign PENetwork_5_io_to_pes_1_out_valid = PE_41_io_data_0_out_valid; // @[pearray.scala 156:36]
  assign PENetwork_5_io_to_pes_1_out_bits = PE_41_io_data_0_out_bits; // @[pearray.scala 156:36]
  assign PENetwork_5_io_to_pes_2_out_valid = PE_42_io_data_0_out_valid; // @[pearray.scala 156:36]
  assign PENetwork_5_io_to_pes_2_out_bits = PE_42_io_data_0_out_bits; // @[pearray.scala 156:36]
  assign PENetwork_5_io_to_pes_3_out_valid = PE_43_io_data_0_out_valid; // @[pearray.scala 156:36]
  assign PENetwork_5_io_to_pes_3_out_bits = PE_43_io_data_0_out_bits; // @[pearray.scala 156:36]
  assign PENetwork_5_io_to_pes_4_out_valid = PE_44_io_data_0_out_valid; // @[pearray.scala 156:36]
  assign PENetwork_5_io_to_pes_4_out_bits = PE_44_io_data_0_out_bits; // @[pearray.scala 156:36]
  assign PENetwork_5_io_to_pes_5_out_valid = PE_45_io_data_0_out_valid; // @[pearray.scala 156:36]
  assign PENetwork_5_io_to_pes_5_out_bits = PE_45_io_data_0_out_bits; // @[pearray.scala 156:36]
  assign PENetwork_5_io_to_pes_6_out_valid = PE_46_io_data_0_out_valid; // @[pearray.scala 156:36]
  assign PENetwork_5_io_to_pes_6_out_bits = PE_46_io_data_0_out_bits; // @[pearray.scala 156:36]
  assign PENetwork_5_io_to_pes_7_out_valid = PE_47_io_data_0_out_valid; // @[pearray.scala 156:36]
  assign PENetwork_5_io_to_pes_7_out_bits = PE_47_io_data_0_out_bits; // @[pearray.scala 156:36]
  assign PENetwork_6_io_to_pes_0_out_valid = PE_48_io_data_0_out_valid; // @[pearray.scala 156:36]
  assign PENetwork_6_io_to_pes_0_out_bits = PE_48_io_data_0_out_bits; // @[pearray.scala 156:36]
  assign PENetwork_6_io_to_pes_1_out_valid = PE_49_io_data_0_out_valid; // @[pearray.scala 156:36]
  assign PENetwork_6_io_to_pes_1_out_bits = PE_49_io_data_0_out_bits; // @[pearray.scala 156:36]
  assign PENetwork_6_io_to_pes_2_out_valid = PE_50_io_data_0_out_valid; // @[pearray.scala 156:36]
  assign PENetwork_6_io_to_pes_2_out_bits = PE_50_io_data_0_out_bits; // @[pearray.scala 156:36]
  assign PENetwork_6_io_to_pes_3_out_valid = PE_51_io_data_0_out_valid; // @[pearray.scala 156:36]
  assign PENetwork_6_io_to_pes_3_out_bits = PE_51_io_data_0_out_bits; // @[pearray.scala 156:36]
  assign PENetwork_6_io_to_pes_4_out_valid = PE_52_io_data_0_out_valid; // @[pearray.scala 156:36]
  assign PENetwork_6_io_to_pes_4_out_bits = PE_52_io_data_0_out_bits; // @[pearray.scala 156:36]
  assign PENetwork_6_io_to_pes_5_out_valid = PE_53_io_data_0_out_valid; // @[pearray.scala 156:36]
  assign PENetwork_6_io_to_pes_5_out_bits = PE_53_io_data_0_out_bits; // @[pearray.scala 156:36]
  assign PENetwork_6_io_to_pes_6_out_valid = PE_54_io_data_0_out_valid; // @[pearray.scala 156:36]
  assign PENetwork_6_io_to_pes_6_out_bits = PE_54_io_data_0_out_bits; // @[pearray.scala 156:36]
  assign PENetwork_6_io_to_pes_7_out_valid = PE_55_io_data_0_out_valid; // @[pearray.scala 156:36]
  assign PENetwork_6_io_to_pes_7_out_bits = PE_55_io_data_0_out_bits; // @[pearray.scala 156:36]
  assign PENetwork_7_io_to_pes_0_out_valid = PE_56_io_data_0_out_valid; // @[pearray.scala 156:36]
  assign PENetwork_7_io_to_pes_0_out_bits = PE_56_io_data_0_out_bits; // @[pearray.scala 156:36]
  assign PENetwork_7_io_to_pes_1_out_valid = PE_57_io_data_0_out_valid; // @[pearray.scala 156:36]
  assign PENetwork_7_io_to_pes_1_out_bits = PE_57_io_data_0_out_bits; // @[pearray.scala 156:36]
  assign PENetwork_7_io_to_pes_2_out_valid = PE_58_io_data_0_out_valid; // @[pearray.scala 156:36]
  assign PENetwork_7_io_to_pes_2_out_bits = PE_58_io_data_0_out_bits; // @[pearray.scala 156:36]
  assign PENetwork_7_io_to_pes_3_out_valid = PE_59_io_data_0_out_valid; // @[pearray.scala 156:36]
  assign PENetwork_7_io_to_pes_3_out_bits = PE_59_io_data_0_out_bits; // @[pearray.scala 156:36]
  assign PENetwork_7_io_to_pes_4_out_valid = PE_60_io_data_0_out_valid; // @[pearray.scala 156:36]
  assign PENetwork_7_io_to_pes_4_out_bits = PE_60_io_data_0_out_bits; // @[pearray.scala 156:36]
  assign PENetwork_7_io_to_pes_5_out_valid = PE_61_io_data_0_out_valid; // @[pearray.scala 156:36]
  assign PENetwork_7_io_to_pes_5_out_bits = PE_61_io_data_0_out_bits; // @[pearray.scala 156:36]
  assign PENetwork_7_io_to_pes_6_out_valid = PE_62_io_data_0_out_valid; // @[pearray.scala 156:36]
  assign PENetwork_7_io_to_pes_6_out_bits = PE_62_io_data_0_out_bits; // @[pearray.scala 156:36]
  assign PENetwork_7_io_to_pes_7_out_valid = PE_63_io_data_0_out_valid; // @[pearray.scala 156:36]
  assign PENetwork_7_io_to_pes_7_out_bits = PE_63_io_data_0_out_bits; // @[pearray.scala 156:36]
  assign PENetwork_8_io_to_pes_0_out_valid = PE_64_io_data_0_out_valid; // @[pearray.scala 156:36]
  assign PENetwork_8_io_to_pes_0_out_bits = PE_64_io_data_0_out_bits; // @[pearray.scala 156:36]
  assign PENetwork_8_io_to_pes_1_out_valid = PE_65_io_data_0_out_valid; // @[pearray.scala 156:36]
  assign PENetwork_8_io_to_pes_1_out_bits = PE_65_io_data_0_out_bits; // @[pearray.scala 156:36]
  assign PENetwork_8_io_to_pes_2_out_valid = PE_66_io_data_0_out_valid; // @[pearray.scala 156:36]
  assign PENetwork_8_io_to_pes_2_out_bits = PE_66_io_data_0_out_bits; // @[pearray.scala 156:36]
  assign PENetwork_8_io_to_pes_3_out_valid = PE_67_io_data_0_out_valid; // @[pearray.scala 156:36]
  assign PENetwork_8_io_to_pes_3_out_bits = PE_67_io_data_0_out_bits; // @[pearray.scala 156:36]
  assign PENetwork_8_io_to_pes_4_out_valid = PE_68_io_data_0_out_valid; // @[pearray.scala 156:36]
  assign PENetwork_8_io_to_pes_4_out_bits = PE_68_io_data_0_out_bits; // @[pearray.scala 156:36]
  assign PENetwork_8_io_to_pes_5_out_valid = PE_69_io_data_0_out_valid; // @[pearray.scala 156:36]
  assign PENetwork_8_io_to_pes_5_out_bits = PE_69_io_data_0_out_bits; // @[pearray.scala 156:36]
  assign PENetwork_8_io_to_pes_6_out_valid = PE_70_io_data_0_out_valid; // @[pearray.scala 156:36]
  assign PENetwork_8_io_to_pes_6_out_bits = PE_70_io_data_0_out_bits; // @[pearray.scala 156:36]
  assign PENetwork_8_io_to_pes_7_out_valid = PE_71_io_data_0_out_valid; // @[pearray.scala 156:36]
  assign PENetwork_8_io_to_pes_7_out_bits = PE_71_io_data_0_out_bits; // @[pearray.scala 156:36]
  assign PENetwork_9_io_to_pes_0_out_valid = PE_72_io_data_0_out_valid; // @[pearray.scala 156:36]
  assign PENetwork_9_io_to_pes_0_out_bits = PE_72_io_data_0_out_bits; // @[pearray.scala 156:36]
  assign PENetwork_9_io_to_pes_1_out_valid = PE_73_io_data_0_out_valid; // @[pearray.scala 156:36]
  assign PENetwork_9_io_to_pes_1_out_bits = PE_73_io_data_0_out_bits; // @[pearray.scala 156:36]
  assign PENetwork_9_io_to_pes_2_out_valid = PE_74_io_data_0_out_valid; // @[pearray.scala 156:36]
  assign PENetwork_9_io_to_pes_2_out_bits = PE_74_io_data_0_out_bits; // @[pearray.scala 156:36]
  assign PENetwork_9_io_to_pes_3_out_valid = PE_75_io_data_0_out_valid; // @[pearray.scala 156:36]
  assign PENetwork_9_io_to_pes_3_out_bits = PE_75_io_data_0_out_bits; // @[pearray.scala 156:36]
  assign PENetwork_9_io_to_pes_4_out_valid = PE_76_io_data_0_out_valid; // @[pearray.scala 156:36]
  assign PENetwork_9_io_to_pes_4_out_bits = PE_76_io_data_0_out_bits; // @[pearray.scala 156:36]
  assign PENetwork_9_io_to_pes_5_out_valid = PE_77_io_data_0_out_valid; // @[pearray.scala 156:36]
  assign PENetwork_9_io_to_pes_5_out_bits = PE_77_io_data_0_out_bits; // @[pearray.scala 156:36]
  assign PENetwork_9_io_to_pes_6_out_valid = PE_78_io_data_0_out_valid; // @[pearray.scala 156:36]
  assign PENetwork_9_io_to_pes_6_out_bits = PE_78_io_data_0_out_bits; // @[pearray.scala 156:36]
  assign PENetwork_9_io_to_pes_7_out_valid = PE_79_io_data_0_out_valid; // @[pearray.scala 156:36]
  assign PENetwork_9_io_to_pes_7_out_bits = PE_79_io_data_0_out_bits; // @[pearray.scala 156:36]
  assign PENetwork_10_io_to_pes_0_out_valid = PE_80_io_data_0_out_valid; // @[pearray.scala 156:36]
  assign PENetwork_10_io_to_pes_0_out_bits = PE_80_io_data_0_out_bits; // @[pearray.scala 156:36]
  assign PENetwork_10_io_to_pes_1_out_valid = PE_81_io_data_0_out_valid; // @[pearray.scala 156:36]
  assign PENetwork_10_io_to_pes_1_out_bits = PE_81_io_data_0_out_bits; // @[pearray.scala 156:36]
  assign PENetwork_10_io_to_pes_2_out_valid = PE_82_io_data_0_out_valid; // @[pearray.scala 156:36]
  assign PENetwork_10_io_to_pes_2_out_bits = PE_82_io_data_0_out_bits; // @[pearray.scala 156:36]
  assign PENetwork_10_io_to_pes_3_out_valid = PE_83_io_data_0_out_valid; // @[pearray.scala 156:36]
  assign PENetwork_10_io_to_pes_3_out_bits = PE_83_io_data_0_out_bits; // @[pearray.scala 156:36]
  assign PENetwork_10_io_to_pes_4_out_valid = PE_84_io_data_0_out_valid; // @[pearray.scala 156:36]
  assign PENetwork_10_io_to_pes_4_out_bits = PE_84_io_data_0_out_bits; // @[pearray.scala 156:36]
  assign PENetwork_10_io_to_pes_5_out_valid = PE_85_io_data_0_out_valid; // @[pearray.scala 156:36]
  assign PENetwork_10_io_to_pes_5_out_bits = PE_85_io_data_0_out_bits; // @[pearray.scala 156:36]
  assign PENetwork_10_io_to_pes_6_out_valid = PE_86_io_data_0_out_valid; // @[pearray.scala 156:36]
  assign PENetwork_10_io_to_pes_6_out_bits = PE_86_io_data_0_out_bits; // @[pearray.scala 156:36]
  assign PENetwork_10_io_to_pes_7_out_valid = PE_87_io_data_0_out_valid; // @[pearray.scala 156:36]
  assign PENetwork_10_io_to_pes_7_out_bits = PE_87_io_data_0_out_bits; // @[pearray.scala 156:36]
  assign PENetwork_11_io_to_pes_0_out_valid = PE_88_io_data_0_out_valid; // @[pearray.scala 156:36]
  assign PENetwork_11_io_to_pes_0_out_bits = PE_88_io_data_0_out_bits; // @[pearray.scala 156:36]
  assign PENetwork_11_io_to_pes_1_out_valid = PE_89_io_data_0_out_valid; // @[pearray.scala 156:36]
  assign PENetwork_11_io_to_pes_1_out_bits = PE_89_io_data_0_out_bits; // @[pearray.scala 156:36]
  assign PENetwork_11_io_to_pes_2_out_valid = PE_90_io_data_0_out_valid; // @[pearray.scala 156:36]
  assign PENetwork_11_io_to_pes_2_out_bits = PE_90_io_data_0_out_bits; // @[pearray.scala 156:36]
  assign PENetwork_11_io_to_pes_3_out_valid = PE_91_io_data_0_out_valid; // @[pearray.scala 156:36]
  assign PENetwork_11_io_to_pes_3_out_bits = PE_91_io_data_0_out_bits; // @[pearray.scala 156:36]
  assign PENetwork_11_io_to_pes_4_out_valid = PE_92_io_data_0_out_valid; // @[pearray.scala 156:36]
  assign PENetwork_11_io_to_pes_4_out_bits = PE_92_io_data_0_out_bits; // @[pearray.scala 156:36]
  assign PENetwork_11_io_to_pes_5_out_valid = PE_93_io_data_0_out_valid; // @[pearray.scala 156:36]
  assign PENetwork_11_io_to_pes_5_out_bits = PE_93_io_data_0_out_bits; // @[pearray.scala 156:36]
  assign PENetwork_11_io_to_pes_6_out_valid = PE_94_io_data_0_out_valid; // @[pearray.scala 156:36]
  assign PENetwork_11_io_to_pes_6_out_bits = PE_94_io_data_0_out_bits; // @[pearray.scala 156:36]
  assign PENetwork_11_io_to_pes_7_out_valid = PE_95_io_data_0_out_valid; // @[pearray.scala 156:36]
  assign PENetwork_11_io_to_pes_7_out_bits = PE_95_io_data_0_out_bits; // @[pearray.scala 156:36]
  assign PENetwork_12_io_to_pes_0_out_valid = PE_96_io_data_0_out_valid; // @[pearray.scala 156:36]
  assign PENetwork_12_io_to_pes_0_out_bits = PE_96_io_data_0_out_bits; // @[pearray.scala 156:36]
  assign PENetwork_12_io_to_pes_1_out_valid = PE_97_io_data_0_out_valid; // @[pearray.scala 156:36]
  assign PENetwork_12_io_to_pes_1_out_bits = PE_97_io_data_0_out_bits; // @[pearray.scala 156:36]
  assign PENetwork_12_io_to_pes_2_out_valid = PE_98_io_data_0_out_valid; // @[pearray.scala 156:36]
  assign PENetwork_12_io_to_pes_2_out_bits = PE_98_io_data_0_out_bits; // @[pearray.scala 156:36]
  assign PENetwork_12_io_to_pes_3_out_valid = PE_99_io_data_0_out_valid; // @[pearray.scala 156:36]
  assign PENetwork_12_io_to_pes_3_out_bits = PE_99_io_data_0_out_bits; // @[pearray.scala 156:36]
  assign PENetwork_12_io_to_pes_4_out_valid = PE_100_io_data_0_out_valid; // @[pearray.scala 156:36]
  assign PENetwork_12_io_to_pes_4_out_bits = PE_100_io_data_0_out_bits; // @[pearray.scala 156:36]
  assign PENetwork_12_io_to_pes_5_out_valid = PE_101_io_data_0_out_valid; // @[pearray.scala 156:36]
  assign PENetwork_12_io_to_pes_5_out_bits = PE_101_io_data_0_out_bits; // @[pearray.scala 156:36]
  assign PENetwork_12_io_to_pes_6_out_valid = PE_102_io_data_0_out_valid; // @[pearray.scala 156:36]
  assign PENetwork_12_io_to_pes_6_out_bits = PE_102_io_data_0_out_bits; // @[pearray.scala 156:36]
  assign PENetwork_12_io_to_pes_7_out_valid = PE_103_io_data_0_out_valid; // @[pearray.scala 156:36]
  assign PENetwork_12_io_to_pes_7_out_bits = PE_103_io_data_0_out_bits; // @[pearray.scala 156:36]
  assign PENetwork_13_io_to_pes_0_out_valid = PE_104_io_data_0_out_valid; // @[pearray.scala 156:36]
  assign PENetwork_13_io_to_pes_0_out_bits = PE_104_io_data_0_out_bits; // @[pearray.scala 156:36]
  assign PENetwork_13_io_to_pes_1_out_valid = PE_105_io_data_0_out_valid; // @[pearray.scala 156:36]
  assign PENetwork_13_io_to_pes_1_out_bits = PE_105_io_data_0_out_bits; // @[pearray.scala 156:36]
  assign PENetwork_13_io_to_pes_2_out_valid = PE_106_io_data_0_out_valid; // @[pearray.scala 156:36]
  assign PENetwork_13_io_to_pes_2_out_bits = PE_106_io_data_0_out_bits; // @[pearray.scala 156:36]
  assign PENetwork_13_io_to_pes_3_out_valid = PE_107_io_data_0_out_valid; // @[pearray.scala 156:36]
  assign PENetwork_13_io_to_pes_3_out_bits = PE_107_io_data_0_out_bits; // @[pearray.scala 156:36]
  assign PENetwork_13_io_to_pes_4_out_valid = PE_108_io_data_0_out_valid; // @[pearray.scala 156:36]
  assign PENetwork_13_io_to_pes_4_out_bits = PE_108_io_data_0_out_bits; // @[pearray.scala 156:36]
  assign PENetwork_13_io_to_pes_5_out_valid = PE_109_io_data_0_out_valid; // @[pearray.scala 156:36]
  assign PENetwork_13_io_to_pes_5_out_bits = PE_109_io_data_0_out_bits; // @[pearray.scala 156:36]
  assign PENetwork_13_io_to_pes_6_out_valid = PE_110_io_data_0_out_valid; // @[pearray.scala 156:36]
  assign PENetwork_13_io_to_pes_6_out_bits = PE_110_io_data_0_out_bits; // @[pearray.scala 156:36]
  assign PENetwork_13_io_to_pes_7_out_valid = PE_111_io_data_0_out_valid; // @[pearray.scala 156:36]
  assign PENetwork_13_io_to_pes_7_out_bits = PE_111_io_data_0_out_bits; // @[pearray.scala 156:36]
  assign PENetwork_14_io_to_pes_0_out_valid = PE_112_io_data_0_out_valid; // @[pearray.scala 156:36]
  assign PENetwork_14_io_to_pes_0_out_bits = PE_112_io_data_0_out_bits; // @[pearray.scala 156:36]
  assign PENetwork_14_io_to_pes_1_out_valid = PE_113_io_data_0_out_valid; // @[pearray.scala 156:36]
  assign PENetwork_14_io_to_pes_1_out_bits = PE_113_io_data_0_out_bits; // @[pearray.scala 156:36]
  assign PENetwork_14_io_to_pes_2_out_valid = PE_114_io_data_0_out_valid; // @[pearray.scala 156:36]
  assign PENetwork_14_io_to_pes_2_out_bits = PE_114_io_data_0_out_bits; // @[pearray.scala 156:36]
  assign PENetwork_14_io_to_pes_3_out_valid = PE_115_io_data_0_out_valid; // @[pearray.scala 156:36]
  assign PENetwork_14_io_to_pes_3_out_bits = PE_115_io_data_0_out_bits; // @[pearray.scala 156:36]
  assign PENetwork_14_io_to_pes_4_out_valid = PE_116_io_data_0_out_valid; // @[pearray.scala 156:36]
  assign PENetwork_14_io_to_pes_4_out_bits = PE_116_io_data_0_out_bits; // @[pearray.scala 156:36]
  assign PENetwork_14_io_to_pes_5_out_valid = PE_117_io_data_0_out_valid; // @[pearray.scala 156:36]
  assign PENetwork_14_io_to_pes_5_out_bits = PE_117_io_data_0_out_bits; // @[pearray.scala 156:36]
  assign PENetwork_14_io_to_pes_6_out_valid = PE_118_io_data_0_out_valid; // @[pearray.scala 156:36]
  assign PENetwork_14_io_to_pes_6_out_bits = PE_118_io_data_0_out_bits; // @[pearray.scala 156:36]
  assign PENetwork_14_io_to_pes_7_out_valid = PE_119_io_data_0_out_valid; // @[pearray.scala 156:36]
  assign PENetwork_14_io_to_pes_7_out_bits = PE_119_io_data_0_out_bits; // @[pearray.scala 156:36]
  assign PENetwork_15_io_to_pes_0_out_valid = PE_120_io_data_0_out_valid; // @[pearray.scala 156:36]
  assign PENetwork_15_io_to_pes_0_out_bits = PE_120_io_data_0_out_bits; // @[pearray.scala 156:36]
  assign PENetwork_15_io_to_pes_1_out_valid = PE_121_io_data_0_out_valid; // @[pearray.scala 156:36]
  assign PENetwork_15_io_to_pes_1_out_bits = PE_121_io_data_0_out_bits; // @[pearray.scala 156:36]
  assign PENetwork_15_io_to_pes_2_out_valid = PE_122_io_data_0_out_valid; // @[pearray.scala 156:36]
  assign PENetwork_15_io_to_pes_2_out_bits = PE_122_io_data_0_out_bits; // @[pearray.scala 156:36]
  assign PENetwork_15_io_to_pes_3_out_valid = PE_123_io_data_0_out_valid; // @[pearray.scala 156:36]
  assign PENetwork_15_io_to_pes_3_out_bits = PE_123_io_data_0_out_bits; // @[pearray.scala 156:36]
  assign PENetwork_15_io_to_pes_4_out_valid = PE_124_io_data_0_out_valid; // @[pearray.scala 156:36]
  assign PENetwork_15_io_to_pes_4_out_bits = PE_124_io_data_0_out_bits; // @[pearray.scala 156:36]
  assign PENetwork_15_io_to_pes_5_out_valid = PE_125_io_data_0_out_valid; // @[pearray.scala 156:36]
  assign PENetwork_15_io_to_pes_5_out_bits = PE_125_io_data_0_out_bits; // @[pearray.scala 156:36]
  assign PENetwork_15_io_to_pes_6_out_valid = PE_126_io_data_0_out_valid; // @[pearray.scala 156:36]
  assign PENetwork_15_io_to_pes_6_out_bits = PE_126_io_data_0_out_bits; // @[pearray.scala 156:36]
  assign PENetwork_15_io_to_pes_7_out_valid = PE_127_io_data_0_out_valid; // @[pearray.scala 156:36]
  assign PENetwork_15_io_to_pes_7_out_bits = PE_127_io_data_0_out_bits; // @[pearray.scala 156:36]
  assign PENetwork_16_io_to_pes_0_out_valid = PE_io_data_1_out_valid; // @[pearray.scala 156:36]
  assign PENetwork_16_io_to_pes_0_out_bits = PE_io_data_1_out_bits; // @[pearray.scala 156:36]
  assign PENetwork_16_io_to_pes_1_out_valid = PE_1_io_data_1_out_valid; // @[pearray.scala 156:36]
  assign PENetwork_16_io_to_pes_1_out_bits = PE_1_io_data_1_out_bits; // @[pearray.scala 156:36]
  assign PENetwork_16_io_to_pes_2_out_valid = PE_2_io_data_1_out_valid; // @[pearray.scala 156:36]
  assign PENetwork_16_io_to_pes_2_out_bits = PE_2_io_data_1_out_bits; // @[pearray.scala 156:36]
  assign PENetwork_16_io_to_pes_3_out_valid = PE_3_io_data_1_out_valid; // @[pearray.scala 156:36]
  assign PENetwork_16_io_to_pes_3_out_bits = PE_3_io_data_1_out_bits; // @[pearray.scala 156:36]
  assign PENetwork_16_io_to_pes_4_out_valid = PE_4_io_data_1_out_valid; // @[pearray.scala 156:36]
  assign PENetwork_16_io_to_pes_4_out_bits = PE_4_io_data_1_out_bits; // @[pearray.scala 156:36]
  assign PENetwork_16_io_to_pes_5_out_valid = PE_5_io_data_1_out_valid; // @[pearray.scala 156:36]
  assign PENetwork_16_io_to_pes_5_out_bits = PE_5_io_data_1_out_bits; // @[pearray.scala 156:36]
  assign PENetwork_16_io_to_pes_6_out_valid = PE_6_io_data_1_out_valid; // @[pearray.scala 156:36]
  assign PENetwork_16_io_to_pes_6_out_bits = PE_6_io_data_1_out_bits; // @[pearray.scala 156:36]
  assign PENetwork_16_io_to_mem_valid = MemController_16_io_rd_data_valid; // @[pearray.scala 239:29]
  assign PENetwork_16_io_to_mem_bits = MemController_16_io_rd_data_bits; // @[pearray.scala 239:29]
  assign PENetwork_17_io_to_pes_0_out_valid = PE_8_io_data_1_out_valid; // @[pearray.scala 156:36]
  assign PENetwork_17_io_to_pes_0_out_bits = PE_8_io_data_1_out_bits; // @[pearray.scala 156:36]
  assign PENetwork_17_io_to_pes_1_out_valid = PE_9_io_data_1_out_valid; // @[pearray.scala 156:36]
  assign PENetwork_17_io_to_pes_1_out_bits = PE_9_io_data_1_out_bits; // @[pearray.scala 156:36]
  assign PENetwork_17_io_to_pes_2_out_valid = PE_10_io_data_1_out_valid; // @[pearray.scala 156:36]
  assign PENetwork_17_io_to_pes_2_out_bits = PE_10_io_data_1_out_bits; // @[pearray.scala 156:36]
  assign PENetwork_17_io_to_pes_3_out_valid = PE_11_io_data_1_out_valid; // @[pearray.scala 156:36]
  assign PENetwork_17_io_to_pes_3_out_bits = PE_11_io_data_1_out_bits; // @[pearray.scala 156:36]
  assign PENetwork_17_io_to_pes_4_out_valid = PE_12_io_data_1_out_valid; // @[pearray.scala 156:36]
  assign PENetwork_17_io_to_pes_4_out_bits = PE_12_io_data_1_out_bits; // @[pearray.scala 156:36]
  assign PENetwork_17_io_to_pes_5_out_valid = PE_13_io_data_1_out_valid; // @[pearray.scala 156:36]
  assign PENetwork_17_io_to_pes_5_out_bits = PE_13_io_data_1_out_bits; // @[pearray.scala 156:36]
  assign PENetwork_17_io_to_pes_6_out_valid = PE_14_io_data_1_out_valid; // @[pearray.scala 156:36]
  assign PENetwork_17_io_to_pes_6_out_bits = PE_14_io_data_1_out_bits; // @[pearray.scala 156:36]
  assign PENetwork_17_io_to_mem_valid = MemController_17_io_rd_data_valid; // @[pearray.scala 239:29]
  assign PENetwork_17_io_to_mem_bits = MemController_17_io_rd_data_bits; // @[pearray.scala 239:29]
  assign PENetwork_18_io_to_pes_0_out_valid = PE_16_io_data_1_out_valid; // @[pearray.scala 156:36]
  assign PENetwork_18_io_to_pes_0_out_bits = PE_16_io_data_1_out_bits; // @[pearray.scala 156:36]
  assign PENetwork_18_io_to_pes_1_out_valid = PE_17_io_data_1_out_valid; // @[pearray.scala 156:36]
  assign PENetwork_18_io_to_pes_1_out_bits = PE_17_io_data_1_out_bits; // @[pearray.scala 156:36]
  assign PENetwork_18_io_to_pes_2_out_valid = PE_18_io_data_1_out_valid; // @[pearray.scala 156:36]
  assign PENetwork_18_io_to_pes_2_out_bits = PE_18_io_data_1_out_bits; // @[pearray.scala 156:36]
  assign PENetwork_18_io_to_pes_3_out_valid = PE_19_io_data_1_out_valid; // @[pearray.scala 156:36]
  assign PENetwork_18_io_to_pes_3_out_bits = PE_19_io_data_1_out_bits; // @[pearray.scala 156:36]
  assign PENetwork_18_io_to_pes_4_out_valid = PE_20_io_data_1_out_valid; // @[pearray.scala 156:36]
  assign PENetwork_18_io_to_pes_4_out_bits = PE_20_io_data_1_out_bits; // @[pearray.scala 156:36]
  assign PENetwork_18_io_to_pes_5_out_valid = PE_21_io_data_1_out_valid; // @[pearray.scala 156:36]
  assign PENetwork_18_io_to_pes_5_out_bits = PE_21_io_data_1_out_bits; // @[pearray.scala 156:36]
  assign PENetwork_18_io_to_pes_6_out_valid = PE_22_io_data_1_out_valid; // @[pearray.scala 156:36]
  assign PENetwork_18_io_to_pes_6_out_bits = PE_22_io_data_1_out_bits; // @[pearray.scala 156:36]
  assign PENetwork_18_io_to_mem_valid = MemController_18_io_rd_data_valid; // @[pearray.scala 239:29]
  assign PENetwork_18_io_to_mem_bits = MemController_18_io_rd_data_bits; // @[pearray.scala 239:29]
  assign PENetwork_19_io_to_pes_0_out_valid = PE_24_io_data_1_out_valid; // @[pearray.scala 156:36]
  assign PENetwork_19_io_to_pes_0_out_bits = PE_24_io_data_1_out_bits; // @[pearray.scala 156:36]
  assign PENetwork_19_io_to_pes_1_out_valid = PE_25_io_data_1_out_valid; // @[pearray.scala 156:36]
  assign PENetwork_19_io_to_pes_1_out_bits = PE_25_io_data_1_out_bits; // @[pearray.scala 156:36]
  assign PENetwork_19_io_to_pes_2_out_valid = PE_26_io_data_1_out_valid; // @[pearray.scala 156:36]
  assign PENetwork_19_io_to_pes_2_out_bits = PE_26_io_data_1_out_bits; // @[pearray.scala 156:36]
  assign PENetwork_19_io_to_pes_3_out_valid = PE_27_io_data_1_out_valid; // @[pearray.scala 156:36]
  assign PENetwork_19_io_to_pes_3_out_bits = PE_27_io_data_1_out_bits; // @[pearray.scala 156:36]
  assign PENetwork_19_io_to_pes_4_out_valid = PE_28_io_data_1_out_valid; // @[pearray.scala 156:36]
  assign PENetwork_19_io_to_pes_4_out_bits = PE_28_io_data_1_out_bits; // @[pearray.scala 156:36]
  assign PENetwork_19_io_to_pes_5_out_valid = PE_29_io_data_1_out_valid; // @[pearray.scala 156:36]
  assign PENetwork_19_io_to_pes_5_out_bits = PE_29_io_data_1_out_bits; // @[pearray.scala 156:36]
  assign PENetwork_19_io_to_pes_6_out_valid = PE_30_io_data_1_out_valid; // @[pearray.scala 156:36]
  assign PENetwork_19_io_to_pes_6_out_bits = PE_30_io_data_1_out_bits; // @[pearray.scala 156:36]
  assign PENetwork_19_io_to_mem_valid = MemController_19_io_rd_data_valid; // @[pearray.scala 239:29]
  assign PENetwork_19_io_to_mem_bits = MemController_19_io_rd_data_bits; // @[pearray.scala 239:29]
  assign PENetwork_20_io_to_pes_0_out_valid = PE_32_io_data_1_out_valid; // @[pearray.scala 156:36]
  assign PENetwork_20_io_to_pes_0_out_bits = PE_32_io_data_1_out_bits; // @[pearray.scala 156:36]
  assign PENetwork_20_io_to_pes_1_out_valid = PE_33_io_data_1_out_valid; // @[pearray.scala 156:36]
  assign PENetwork_20_io_to_pes_1_out_bits = PE_33_io_data_1_out_bits; // @[pearray.scala 156:36]
  assign PENetwork_20_io_to_pes_2_out_valid = PE_34_io_data_1_out_valid; // @[pearray.scala 156:36]
  assign PENetwork_20_io_to_pes_2_out_bits = PE_34_io_data_1_out_bits; // @[pearray.scala 156:36]
  assign PENetwork_20_io_to_pes_3_out_valid = PE_35_io_data_1_out_valid; // @[pearray.scala 156:36]
  assign PENetwork_20_io_to_pes_3_out_bits = PE_35_io_data_1_out_bits; // @[pearray.scala 156:36]
  assign PENetwork_20_io_to_pes_4_out_valid = PE_36_io_data_1_out_valid; // @[pearray.scala 156:36]
  assign PENetwork_20_io_to_pes_4_out_bits = PE_36_io_data_1_out_bits; // @[pearray.scala 156:36]
  assign PENetwork_20_io_to_pes_5_out_valid = PE_37_io_data_1_out_valid; // @[pearray.scala 156:36]
  assign PENetwork_20_io_to_pes_5_out_bits = PE_37_io_data_1_out_bits; // @[pearray.scala 156:36]
  assign PENetwork_20_io_to_pes_6_out_valid = PE_38_io_data_1_out_valid; // @[pearray.scala 156:36]
  assign PENetwork_20_io_to_pes_6_out_bits = PE_38_io_data_1_out_bits; // @[pearray.scala 156:36]
  assign PENetwork_20_io_to_mem_valid = MemController_20_io_rd_data_valid; // @[pearray.scala 239:29]
  assign PENetwork_20_io_to_mem_bits = MemController_20_io_rd_data_bits; // @[pearray.scala 239:29]
  assign PENetwork_21_io_to_pes_0_out_valid = PE_40_io_data_1_out_valid; // @[pearray.scala 156:36]
  assign PENetwork_21_io_to_pes_0_out_bits = PE_40_io_data_1_out_bits; // @[pearray.scala 156:36]
  assign PENetwork_21_io_to_pes_1_out_valid = PE_41_io_data_1_out_valid; // @[pearray.scala 156:36]
  assign PENetwork_21_io_to_pes_1_out_bits = PE_41_io_data_1_out_bits; // @[pearray.scala 156:36]
  assign PENetwork_21_io_to_pes_2_out_valid = PE_42_io_data_1_out_valid; // @[pearray.scala 156:36]
  assign PENetwork_21_io_to_pes_2_out_bits = PE_42_io_data_1_out_bits; // @[pearray.scala 156:36]
  assign PENetwork_21_io_to_pes_3_out_valid = PE_43_io_data_1_out_valid; // @[pearray.scala 156:36]
  assign PENetwork_21_io_to_pes_3_out_bits = PE_43_io_data_1_out_bits; // @[pearray.scala 156:36]
  assign PENetwork_21_io_to_pes_4_out_valid = PE_44_io_data_1_out_valid; // @[pearray.scala 156:36]
  assign PENetwork_21_io_to_pes_4_out_bits = PE_44_io_data_1_out_bits; // @[pearray.scala 156:36]
  assign PENetwork_21_io_to_pes_5_out_valid = PE_45_io_data_1_out_valid; // @[pearray.scala 156:36]
  assign PENetwork_21_io_to_pes_5_out_bits = PE_45_io_data_1_out_bits; // @[pearray.scala 156:36]
  assign PENetwork_21_io_to_pes_6_out_valid = PE_46_io_data_1_out_valid; // @[pearray.scala 156:36]
  assign PENetwork_21_io_to_pes_6_out_bits = PE_46_io_data_1_out_bits; // @[pearray.scala 156:36]
  assign PENetwork_21_io_to_mem_valid = MemController_21_io_rd_data_valid; // @[pearray.scala 239:29]
  assign PENetwork_21_io_to_mem_bits = MemController_21_io_rd_data_bits; // @[pearray.scala 239:29]
  assign PENetwork_22_io_to_pes_0_out_valid = PE_48_io_data_1_out_valid; // @[pearray.scala 156:36]
  assign PENetwork_22_io_to_pes_0_out_bits = PE_48_io_data_1_out_bits; // @[pearray.scala 156:36]
  assign PENetwork_22_io_to_pes_1_out_valid = PE_49_io_data_1_out_valid; // @[pearray.scala 156:36]
  assign PENetwork_22_io_to_pes_1_out_bits = PE_49_io_data_1_out_bits; // @[pearray.scala 156:36]
  assign PENetwork_22_io_to_pes_2_out_valid = PE_50_io_data_1_out_valid; // @[pearray.scala 156:36]
  assign PENetwork_22_io_to_pes_2_out_bits = PE_50_io_data_1_out_bits; // @[pearray.scala 156:36]
  assign PENetwork_22_io_to_pes_3_out_valid = PE_51_io_data_1_out_valid; // @[pearray.scala 156:36]
  assign PENetwork_22_io_to_pes_3_out_bits = PE_51_io_data_1_out_bits; // @[pearray.scala 156:36]
  assign PENetwork_22_io_to_pes_4_out_valid = PE_52_io_data_1_out_valid; // @[pearray.scala 156:36]
  assign PENetwork_22_io_to_pes_4_out_bits = PE_52_io_data_1_out_bits; // @[pearray.scala 156:36]
  assign PENetwork_22_io_to_pes_5_out_valid = PE_53_io_data_1_out_valid; // @[pearray.scala 156:36]
  assign PENetwork_22_io_to_pes_5_out_bits = PE_53_io_data_1_out_bits; // @[pearray.scala 156:36]
  assign PENetwork_22_io_to_pes_6_out_valid = PE_54_io_data_1_out_valid; // @[pearray.scala 156:36]
  assign PENetwork_22_io_to_pes_6_out_bits = PE_54_io_data_1_out_bits; // @[pearray.scala 156:36]
  assign PENetwork_22_io_to_mem_valid = MemController_22_io_rd_data_valid; // @[pearray.scala 239:29]
  assign PENetwork_22_io_to_mem_bits = MemController_22_io_rd_data_bits; // @[pearray.scala 239:29]
  assign PENetwork_23_io_to_pes_0_out_valid = PE_56_io_data_1_out_valid; // @[pearray.scala 156:36]
  assign PENetwork_23_io_to_pes_0_out_bits = PE_56_io_data_1_out_bits; // @[pearray.scala 156:36]
  assign PENetwork_23_io_to_pes_1_out_valid = PE_57_io_data_1_out_valid; // @[pearray.scala 156:36]
  assign PENetwork_23_io_to_pes_1_out_bits = PE_57_io_data_1_out_bits; // @[pearray.scala 156:36]
  assign PENetwork_23_io_to_pes_2_out_valid = PE_58_io_data_1_out_valid; // @[pearray.scala 156:36]
  assign PENetwork_23_io_to_pes_2_out_bits = PE_58_io_data_1_out_bits; // @[pearray.scala 156:36]
  assign PENetwork_23_io_to_pes_3_out_valid = PE_59_io_data_1_out_valid; // @[pearray.scala 156:36]
  assign PENetwork_23_io_to_pes_3_out_bits = PE_59_io_data_1_out_bits; // @[pearray.scala 156:36]
  assign PENetwork_23_io_to_pes_4_out_valid = PE_60_io_data_1_out_valid; // @[pearray.scala 156:36]
  assign PENetwork_23_io_to_pes_4_out_bits = PE_60_io_data_1_out_bits; // @[pearray.scala 156:36]
  assign PENetwork_23_io_to_pes_5_out_valid = PE_61_io_data_1_out_valid; // @[pearray.scala 156:36]
  assign PENetwork_23_io_to_pes_5_out_bits = PE_61_io_data_1_out_bits; // @[pearray.scala 156:36]
  assign PENetwork_23_io_to_pes_6_out_valid = PE_62_io_data_1_out_valid; // @[pearray.scala 156:36]
  assign PENetwork_23_io_to_pes_6_out_bits = PE_62_io_data_1_out_bits; // @[pearray.scala 156:36]
  assign PENetwork_23_io_to_mem_valid = MemController_23_io_rd_data_valid; // @[pearray.scala 239:29]
  assign PENetwork_23_io_to_mem_bits = MemController_23_io_rd_data_bits; // @[pearray.scala 239:29]
  assign PENetwork_24_io_to_pes_0_out_valid = PE_64_io_data_1_out_valid; // @[pearray.scala 156:36]
  assign PENetwork_24_io_to_pes_0_out_bits = PE_64_io_data_1_out_bits; // @[pearray.scala 156:36]
  assign PENetwork_24_io_to_pes_1_out_valid = PE_65_io_data_1_out_valid; // @[pearray.scala 156:36]
  assign PENetwork_24_io_to_pes_1_out_bits = PE_65_io_data_1_out_bits; // @[pearray.scala 156:36]
  assign PENetwork_24_io_to_pes_2_out_valid = PE_66_io_data_1_out_valid; // @[pearray.scala 156:36]
  assign PENetwork_24_io_to_pes_2_out_bits = PE_66_io_data_1_out_bits; // @[pearray.scala 156:36]
  assign PENetwork_24_io_to_pes_3_out_valid = PE_67_io_data_1_out_valid; // @[pearray.scala 156:36]
  assign PENetwork_24_io_to_pes_3_out_bits = PE_67_io_data_1_out_bits; // @[pearray.scala 156:36]
  assign PENetwork_24_io_to_pes_4_out_valid = PE_68_io_data_1_out_valid; // @[pearray.scala 156:36]
  assign PENetwork_24_io_to_pes_4_out_bits = PE_68_io_data_1_out_bits; // @[pearray.scala 156:36]
  assign PENetwork_24_io_to_pes_5_out_valid = PE_69_io_data_1_out_valid; // @[pearray.scala 156:36]
  assign PENetwork_24_io_to_pes_5_out_bits = PE_69_io_data_1_out_bits; // @[pearray.scala 156:36]
  assign PENetwork_24_io_to_pes_6_out_valid = PE_70_io_data_1_out_valid; // @[pearray.scala 156:36]
  assign PENetwork_24_io_to_pes_6_out_bits = PE_70_io_data_1_out_bits; // @[pearray.scala 156:36]
  assign PENetwork_24_io_to_mem_valid = MemController_24_io_rd_data_valid; // @[pearray.scala 239:29]
  assign PENetwork_24_io_to_mem_bits = MemController_24_io_rd_data_bits; // @[pearray.scala 239:29]
  assign PENetwork_25_io_to_pes_0_out_valid = PE_72_io_data_1_out_valid; // @[pearray.scala 156:36]
  assign PENetwork_25_io_to_pes_0_out_bits = PE_72_io_data_1_out_bits; // @[pearray.scala 156:36]
  assign PENetwork_25_io_to_pes_1_out_valid = PE_73_io_data_1_out_valid; // @[pearray.scala 156:36]
  assign PENetwork_25_io_to_pes_1_out_bits = PE_73_io_data_1_out_bits; // @[pearray.scala 156:36]
  assign PENetwork_25_io_to_pes_2_out_valid = PE_74_io_data_1_out_valid; // @[pearray.scala 156:36]
  assign PENetwork_25_io_to_pes_2_out_bits = PE_74_io_data_1_out_bits; // @[pearray.scala 156:36]
  assign PENetwork_25_io_to_pes_3_out_valid = PE_75_io_data_1_out_valid; // @[pearray.scala 156:36]
  assign PENetwork_25_io_to_pes_3_out_bits = PE_75_io_data_1_out_bits; // @[pearray.scala 156:36]
  assign PENetwork_25_io_to_pes_4_out_valid = PE_76_io_data_1_out_valid; // @[pearray.scala 156:36]
  assign PENetwork_25_io_to_pes_4_out_bits = PE_76_io_data_1_out_bits; // @[pearray.scala 156:36]
  assign PENetwork_25_io_to_pes_5_out_valid = PE_77_io_data_1_out_valid; // @[pearray.scala 156:36]
  assign PENetwork_25_io_to_pes_5_out_bits = PE_77_io_data_1_out_bits; // @[pearray.scala 156:36]
  assign PENetwork_25_io_to_pes_6_out_valid = PE_78_io_data_1_out_valid; // @[pearray.scala 156:36]
  assign PENetwork_25_io_to_pes_6_out_bits = PE_78_io_data_1_out_bits; // @[pearray.scala 156:36]
  assign PENetwork_25_io_to_mem_valid = MemController_25_io_rd_data_valid; // @[pearray.scala 239:29]
  assign PENetwork_25_io_to_mem_bits = MemController_25_io_rd_data_bits; // @[pearray.scala 239:29]
  assign PENetwork_26_io_to_pes_0_out_valid = PE_80_io_data_1_out_valid; // @[pearray.scala 156:36]
  assign PENetwork_26_io_to_pes_0_out_bits = PE_80_io_data_1_out_bits; // @[pearray.scala 156:36]
  assign PENetwork_26_io_to_pes_1_out_valid = PE_81_io_data_1_out_valid; // @[pearray.scala 156:36]
  assign PENetwork_26_io_to_pes_1_out_bits = PE_81_io_data_1_out_bits; // @[pearray.scala 156:36]
  assign PENetwork_26_io_to_pes_2_out_valid = PE_82_io_data_1_out_valid; // @[pearray.scala 156:36]
  assign PENetwork_26_io_to_pes_2_out_bits = PE_82_io_data_1_out_bits; // @[pearray.scala 156:36]
  assign PENetwork_26_io_to_pes_3_out_valid = PE_83_io_data_1_out_valid; // @[pearray.scala 156:36]
  assign PENetwork_26_io_to_pes_3_out_bits = PE_83_io_data_1_out_bits; // @[pearray.scala 156:36]
  assign PENetwork_26_io_to_pes_4_out_valid = PE_84_io_data_1_out_valid; // @[pearray.scala 156:36]
  assign PENetwork_26_io_to_pes_4_out_bits = PE_84_io_data_1_out_bits; // @[pearray.scala 156:36]
  assign PENetwork_26_io_to_pes_5_out_valid = PE_85_io_data_1_out_valid; // @[pearray.scala 156:36]
  assign PENetwork_26_io_to_pes_5_out_bits = PE_85_io_data_1_out_bits; // @[pearray.scala 156:36]
  assign PENetwork_26_io_to_pes_6_out_valid = PE_86_io_data_1_out_valid; // @[pearray.scala 156:36]
  assign PENetwork_26_io_to_pes_6_out_bits = PE_86_io_data_1_out_bits; // @[pearray.scala 156:36]
  assign PENetwork_26_io_to_mem_valid = MemController_26_io_rd_data_valid; // @[pearray.scala 239:29]
  assign PENetwork_26_io_to_mem_bits = MemController_26_io_rd_data_bits; // @[pearray.scala 239:29]
  assign PENetwork_27_io_to_pes_0_out_valid = PE_88_io_data_1_out_valid; // @[pearray.scala 156:36]
  assign PENetwork_27_io_to_pes_0_out_bits = PE_88_io_data_1_out_bits; // @[pearray.scala 156:36]
  assign PENetwork_27_io_to_pes_1_out_valid = PE_89_io_data_1_out_valid; // @[pearray.scala 156:36]
  assign PENetwork_27_io_to_pes_1_out_bits = PE_89_io_data_1_out_bits; // @[pearray.scala 156:36]
  assign PENetwork_27_io_to_pes_2_out_valid = PE_90_io_data_1_out_valid; // @[pearray.scala 156:36]
  assign PENetwork_27_io_to_pes_2_out_bits = PE_90_io_data_1_out_bits; // @[pearray.scala 156:36]
  assign PENetwork_27_io_to_pes_3_out_valid = PE_91_io_data_1_out_valid; // @[pearray.scala 156:36]
  assign PENetwork_27_io_to_pes_3_out_bits = PE_91_io_data_1_out_bits; // @[pearray.scala 156:36]
  assign PENetwork_27_io_to_pes_4_out_valid = PE_92_io_data_1_out_valid; // @[pearray.scala 156:36]
  assign PENetwork_27_io_to_pes_4_out_bits = PE_92_io_data_1_out_bits; // @[pearray.scala 156:36]
  assign PENetwork_27_io_to_pes_5_out_valid = PE_93_io_data_1_out_valid; // @[pearray.scala 156:36]
  assign PENetwork_27_io_to_pes_5_out_bits = PE_93_io_data_1_out_bits; // @[pearray.scala 156:36]
  assign PENetwork_27_io_to_pes_6_out_valid = PE_94_io_data_1_out_valid; // @[pearray.scala 156:36]
  assign PENetwork_27_io_to_pes_6_out_bits = PE_94_io_data_1_out_bits; // @[pearray.scala 156:36]
  assign PENetwork_27_io_to_mem_valid = MemController_27_io_rd_data_valid; // @[pearray.scala 239:29]
  assign PENetwork_27_io_to_mem_bits = MemController_27_io_rd_data_bits; // @[pearray.scala 239:29]
  assign PENetwork_28_io_to_pes_0_out_valid = PE_96_io_data_1_out_valid; // @[pearray.scala 156:36]
  assign PENetwork_28_io_to_pes_0_out_bits = PE_96_io_data_1_out_bits; // @[pearray.scala 156:36]
  assign PENetwork_28_io_to_pes_1_out_valid = PE_97_io_data_1_out_valid; // @[pearray.scala 156:36]
  assign PENetwork_28_io_to_pes_1_out_bits = PE_97_io_data_1_out_bits; // @[pearray.scala 156:36]
  assign PENetwork_28_io_to_pes_2_out_valid = PE_98_io_data_1_out_valid; // @[pearray.scala 156:36]
  assign PENetwork_28_io_to_pes_2_out_bits = PE_98_io_data_1_out_bits; // @[pearray.scala 156:36]
  assign PENetwork_28_io_to_pes_3_out_valid = PE_99_io_data_1_out_valid; // @[pearray.scala 156:36]
  assign PENetwork_28_io_to_pes_3_out_bits = PE_99_io_data_1_out_bits; // @[pearray.scala 156:36]
  assign PENetwork_28_io_to_pes_4_out_valid = PE_100_io_data_1_out_valid; // @[pearray.scala 156:36]
  assign PENetwork_28_io_to_pes_4_out_bits = PE_100_io_data_1_out_bits; // @[pearray.scala 156:36]
  assign PENetwork_28_io_to_pes_5_out_valid = PE_101_io_data_1_out_valid; // @[pearray.scala 156:36]
  assign PENetwork_28_io_to_pes_5_out_bits = PE_101_io_data_1_out_bits; // @[pearray.scala 156:36]
  assign PENetwork_28_io_to_pes_6_out_valid = PE_102_io_data_1_out_valid; // @[pearray.scala 156:36]
  assign PENetwork_28_io_to_pes_6_out_bits = PE_102_io_data_1_out_bits; // @[pearray.scala 156:36]
  assign PENetwork_28_io_to_mem_valid = MemController_28_io_rd_data_valid; // @[pearray.scala 239:29]
  assign PENetwork_28_io_to_mem_bits = MemController_28_io_rd_data_bits; // @[pearray.scala 239:29]
  assign PENetwork_29_io_to_pes_0_out_valid = PE_104_io_data_1_out_valid; // @[pearray.scala 156:36]
  assign PENetwork_29_io_to_pes_0_out_bits = PE_104_io_data_1_out_bits; // @[pearray.scala 156:36]
  assign PENetwork_29_io_to_pes_1_out_valid = PE_105_io_data_1_out_valid; // @[pearray.scala 156:36]
  assign PENetwork_29_io_to_pes_1_out_bits = PE_105_io_data_1_out_bits; // @[pearray.scala 156:36]
  assign PENetwork_29_io_to_pes_2_out_valid = PE_106_io_data_1_out_valid; // @[pearray.scala 156:36]
  assign PENetwork_29_io_to_pes_2_out_bits = PE_106_io_data_1_out_bits; // @[pearray.scala 156:36]
  assign PENetwork_29_io_to_pes_3_out_valid = PE_107_io_data_1_out_valid; // @[pearray.scala 156:36]
  assign PENetwork_29_io_to_pes_3_out_bits = PE_107_io_data_1_out_bits; // @[pearray.scala 156:36]
  assign PENetwork_29_io_to_pes_4_out_valid = PE_108_io_data_1_out_valid; // @[pearray.scala 156:36]
  assign PENetwork_29_io_to_pes_4_out_bits = PE_108_io_data_1_out_bits; // @[pearray.scala 156:36]
  assign PENetwork_29_io_to_pes_5_out_valid = PE_109_io_data_1_out_valid; // @[pearray.scala 156:36]
  assign PENetwork_29_io_to_pes_5_out_bits = PE_109_io_data_1_out_bits; // @[pearray.scala 156:36]
  assign PENetwork_29_io_to_pes_6_out_valid = PE_110_io_data_1_out_valid; // @[pearray.scala 156:36]
  assign PENetwork_29_io_to_pes_6_out_bits = PE_110_io_data_1_out_bits; // @[pearray.scala 156:36]
  assign PENetwork_29_io_to_mem_valid = MemController_29_io_rd_data_valid; // @[pearray.scala 239:29]
  assign PENetwork_29_io_to_mem_bits = MemController_29_io_rd_data_bits; // @[pearray.scala 239:29]
  assign PENetwork_30_io_to_pes_0_out_valid = PE_112_io_data_1_out_valid; // @[pearray.scala 156:36]
  assign PENetwork_30_io_to_pes_0_out_bits = PE_112_io_data_1_out_bits; // @[pearray.scala 156:36]
  assign PENetwork_30_io_to_pes_1_out_valid = PE_113_io_data_1_out_valid; // @[pearray.scala 156:36]
  assign PENetwork_30_io_to_pes_1_out_bits = PE_113_io_data_1_out_bits; // @[pearray.scala 156:36]
  assign PENetwork_30_io_to_pes_2_out_valid = PE_114_io_data_1_out_valid; // @[pearray.scala 156:36]
  assign PENetwork_30_io_to_pes_2_out_bits = PE_114_io_data_1_out_bits; // @[pearray.scala 156:36]
  assign PENetwork_30_io_to_pes_3_out_valid = PE_115_io_data_1_out_valid; // @[pearray.scala 156:36]
  assign PENetwork_30_io_to_pes_3_out_bits = PE_115_io_data_1_out_bits; // @[pearray.scala 156:36]
  assign PENetwork_30_io_to_pes_4_out_valid = PE_116_io_data_1_out_valid; // @[pearray.scala 156:36]
  assign PENetwork_30_io_to_pes_4_out_bits = PE_116_io_data_1_out_bits; // @[pearray.scala 156:36]
  assign PENetwork_30_io_to_pes_5_out_valid = PE_117_io_data_1_out_valid; // @[pearray.scala 156:36]
  assign PENetwork_30_io_to_pes_5_out_bits = PE_117_io_data_1_out_bits; // @[pearray.scala 156:36]
  assign PENetwork_30_io_to_pes_6_out_valid = PE_118_io_data_1_out_valid; // @[pearray.scala 156:36]
  assign PENetwork_30_io_to_pes_6_out_bits = PE_118_io_data_1_out_bits; // @[pearray.scala 156:36]
  assign PENetwork_30_io_to_mem_valid = MemController_30_io_rd_data_valid; // @[pearray.scala 239:29]
  assign PENetwork_30_io_to_mem_bits = MemController_30_io_rd_data_bits; // @[pearray.scala 239:29]
  assign PENetwork_31_io_to_pes_0_out_valid = PE_120_io_data_1_out_valid; // @[pearray.scala 156:36]
  assign PENetwork_31_io_to_pes_0_out_bits = PE_120_io_data_1_out_bits; // @[pearray.scala 156:36]
  assign PENetwork_31_io_to_pes_1_out_valid = PE_121_io_data_1_out_valid; // @[pearray.scala 156:36]
  assign PENetwork_31_io_to_pes_1_out_bits = PE_121_io_data_1_out_bits; // @[pearray.scala 156:36]
  assign PENetwork_31_io_to_pes_2_out_valid = PE_122_io_data_1_out_valid; // @[pearray.scala 156:36]
  assign PENetwork_31_io_to_pes_2_out_bits = PE_122_io_data_1_out_bits; // @[pearray.scala 156:36]
  assign PENetwork_31_io_to_pes_3_out_valid = PE_123_io_data_1_out_valid; // @[pearray.scala 156:36]
  assign PENetwork_31_io_to_pes_3_out_bits = PE_123_io_data_1_out_bits; // @[pearray.scala 156:36]
  assign PENetwork_31_io_to_pes_4_out_valid = PE_124_io_data_1_out_valid; // @[pearray.scala 156:36]
  assign PENetwork_31_io_to_pes_4_out_bits = PE_124_io_data_1_out_bits; // @[pearray.scala 156:36]
  assign PENetwork_31_io_to_pes_5_out_valid = PE_125_io_data_1_out_valid; // @[pearray.scala 156:36]
  assign PENetwork_31_io_to_pes_5_out_bits = PE_125_io_data_1_out_bits; // @[pearray.scala 156:36]
  assign PENetwork_31_io_to_pes_6_out_valid = PE_126_io_data_1_out_valid; // @[pearray.scala 156:36]
  assign PENetwork_31_io_to_pes_6_out_bits = PE_126_io_data_1_out_bits; // @[pearray.scala 156:36]
  assign PENetwork_31_io_to_mem_valid = MemController_31_io_rd_data_valid; // @[pearray.scala 239:29]
  assign PENetwork_31_io_to_mem_bits = MemController_31_io_rd_data_bits; // @[pearray.scala 239:29]
  assign PENetwork_32_io_to_pes_0_out_bits = PE_io_data_2_out_bits; // @[pearray.scala 156:36]
  assign PENetwork_32_io_to_pes_1_out_bits = PE_8_io_data_2_out_bits; // @[pearray.scala 156:36]
  assign PENetwork_32_io_to_pes_2_out_bits = PE_16_io_data_2_out_bits; // @[pearray.scala 156:36]
  assign PENetwork_32_io_to_pes_3_out_bits = PE_24_io_data_2_out_bits; // @[pearray.scala 156:36]
  assign PENetwork_32_io_to_pes_4_out_bits = PE_32_io_data_2_out_bits; // @[pearray.scala 156:36]
  assign PENetwork_32_io_to_pes_5_out_bits = PE_40_io_data_2_out_bits; // @[pearray.scala 156:36]
  assign PENetwork_32_io_to_pes_6_out_bits = PE_48_io_data_2_out_bits; // @[pearray.scala 156:36]
  assign PENetwork_32_io_to_pes_7_out_bits = PE_56_io_data_2_out_bits; // @[pearray.scala 156:36]
  assign PENetwork_32_io_to_pes_8_out_bits = PE_64_io_data_2_out_bits; // @[pearray.scala 156:36]
  assign PENetwork_32_io_to_pes_9_out_bits = PE_72_io_data_2_out_bits; // @[pearray.scala 156:36]
  assign PENetwork_32_io_to_pes_10_out_bits = PE_80_io_data_2_out_bits; // @[pearray.scala 156:36]
  assign PENetwork_32_io_to_pes_11_out_bits = PE_88_io_data_2_out_bits; // @[pearray.scala 156:36]
  assign PENetwork_32_io_to_pes_12_out_bits = PE_96_io_data_2_out_bits; // @[pearray.scala 156:36]
  assign PENetwork_32_io_to_pes_13_out_bits = PE_104_io_data_2_out_bits; // @[pearray.scala 156:36]
  assign PENetwork_32_io_to_pes_14_out_bits = PE_112_io_data_2_out_bits; // @[pearray.scala 156:36]
  assign PENetwork_32_io_to_mem_bits = MemController_32_io_rd_data_bits; // @[pearray.scala 239:29]
  assign PENetwork_33_io_to_pes_0_out_bits = PE_1_io_data_2_out_bits; // @[pearray.scala 156:36]
  assign PENetwork_33_io_to_pes_1_out_bits = PE_9_io_data_2_out_bits; // @[pearray.scala 156:36]
  assign PENetwork_33_io_to_pes_2_out_bits = PE_17_io_data_2_out_bits; // @[pearray.scala 156:36]
  assign PENetwork_33_io_to_pes_3_out_bits = PE_25_io_data_2_out_bits; // @[pearray.scala 156:36]
  assign PENetwork_33_io_to_pes_4_out_bits = PE_33_io_data_2_out_bits; // @[pearray.scala 156:36]
  assign PENetwork_33_io_to_pes_5_out_bits = PE_41_io_data_2_out_bits; // @[pearray.scala 156:36]
  assign PENetwork_33_io_to_pes_6_out_bits = PE_49_io_data_2_out_bits; // @[pearray.scala 156:36]
  assign PENetwork_33_io_to_pes_7_out_bits = PE_57_io_data_2_out_bits; // @[pearray.scala 156:36]
  assign PENetwork_33_io_to_pes_8_out_bits = PE_65_io_data_2_out_bits; // @[pearray.scala 156:36]
  assign PENetwork_33_io_to_pes_9_out_bits = PE_73_io_data_2_out_bits; // @[pearray.scala 156:36]
  assign PENetwork_33_io_to_pes_10_out_bits = PE_81_io_data_2_out_bits; // @[pearray.scala 156:36]
  assign PENetwork_33_io_to_pes_11_out_bits = PE_89_io_data_2_out_bits; // @[pearray.scala 156:36]
  assign PENetwork_33_io_to_pes_12_out_bits = PE_97_io_data_2_out_bits; // @[pearray.scala 156:36]
  assign PENetwork_33_io_to_pes_13_out_bits = PE_105_io_data_2_out_bits; // @[pearray.scala 156:36]
  assign PENetwork_33_io_to_pes_14_out_bits = PE_113_io_data_2_out_bits; // @[pearray.scala 156:36]
  assign PENetwork_33_io_to_mem_bits = MemController_33_io_rd_data_bits; // @[pearray.scala 239:29]
  assign PENetwork_34_io_to_pes_0_out_bits = PE_2_io_data_2_out_bits; // @[pearray.scala 156:36]
  assign PENetwork_34_io_to_pes_1_out_bits = PE_10_io_data_2_out_bits; // @[pearray.scala 156:36]
  assign PENetwork_34_io_to_pes_2_out_bits = PE_18_io_data_2_out_bits; // @[pearray.scala 156:36]
  assign PENetwork_34_io_to_pes_3_out_bits = PE_26_io_data_2_out_bits; // @[pearray.scala 156:36]
  assign PENetwork_34_io_to_pes_4_out_bits = PE_34_io_data_2_out_bits; // @[pearray.scala 156:36]
  assign PENetwork_34_io_to_pes_5_out_bits = PE_42_io_data_2_out_bits; // @[pearray.scala 156:36]
  assign PENetwork_34_io_to_pes_6_out_bits = PE_50_io_data_2_out_bits; // @[pearray.scala 156:36]
  assign PENetwork_34_io_to_pes_7_out_bits = PE_58_io_data_2_out_bits; // @[pearray.scala 156:36]
  assign PENetwork_34_io_to_pes_8_out_bits = PE_66_io_data_2_out_bits; // @[pearray.scala 156:36]
  assign PENetwork_34_io_to_pes_9_out_bits = PE_74_io_data_2_out_bits; // @[pearray.scala 156:36]
  assign PENetwork_34_io_to_pes_10_out_bits = PE_82_io_data_2_out_bits; // @[pearray.scala 156:36]
  assign PENetwork_34_io_to_pes_11_out_bits = PE_90_io_data_2_out_bits; // @[pearray.scala 156:36]
  assign PENetwork_34_io_to_pes_12_out_bits = PE_98_io_data_2_out_bits; // @[pearray.scala 156:36]
  assign PENetwork_34_io_to_pes_13_out_bits = PE_106_io_data_2_out_bits; // @[pearray.scala 156:36]
  assign PENetwork_34_io_to_pes_14_out_bits = PE_114_io_data_2_out_bits; // @[pearray.scala 156:36]
  assign PENetwork_34_io_to_mem_bits = MemController_34_io_rd_data_bits; // @[pearray.scala 239:29]
  assign PENetwork_35_io_to_pes_0_out_bits = PE_3_io_data_2_out_bits; // @[pearray.scala 156:36]
  assign PENetwork_35_io_to_pes_1_out_bits = PE_11_io_data_2_out_bits; // @[pearray.scala 156:36]
  assign PENetwork_35_io_to_pes_2_out_bits = PE_19_io_data_2_out_bits; // @[pearray.scala 156:36]
  assign PENetwork_35_io_to_pes_3_out_bits = PE_27_io_data_2_out_bits; // @[pearray.scala 156:36]
  assign PENetwork_35_io_to_pes_4_out_bits = PE_35_io_data_2_out_bits; // @[pearray.scala 156:36]
  assign PENetwork_35_io_to_pes_5_out_bits = PE_43_io_data_2_out_bits; // @[pearray.scala 156:36]
  assign PENetwork_35_io_to_pes_6_out_bits = PE_51_io_data_2_out_bits; // @[pearray.scala 156:36]
  assign PENetwork_35_io_to_pes_7_out_bits = PE_59_io_data_2_out_bits; // @[pearray.scala 156:36]
  assign PENetwork_35_io_to_pes_8_out_bits = PE_67_io_data_2_out_bits; // @[pearray.scala 156:36]
  assign PENetwork_35_io_to_pes_9_out_bits = PE_75_io_data_2_out_bits; // @[pearray.scala 156:36]
  assign PENetwork_35_io_to_pes_10_out_bits = PE_83_io_data_2_out_bits; // @[pearray.scala 156:36]
  assign PENetwork_35_io_to_pes_11_out_bits = PE_91_io_data_2_out_bits; // @[pearray.scala 156:36]
  assign PENetwork_35_io_to_pes_12_out_bits = PE_99_io_data_2_out_bits; // @[pearray.scala 156:36]
  assign PENetwork_35_io_to_pes_13_out_bits = PE_107_io_data_2_out_bits; // @[pearray.scala 156:36]
  assign PENetwork_35_io_to_pes_14_out_bits = PE_115_io_data_2_out_bits; // @[pearray.scala 156:36]
  assign PENetwork_35_io_to_mem_bits = MemController_35_io_rd_data_bits; // @[pearray.scala 239:29]
  assign PENetwork_36_io_to_pes_0_out_bits = PE_4_io_data_2_out_bits; // @[pearray.scala 156:36]
  assign PENetwork_36_io_to_pes_1_out_bits = PE_12_io_data_2_out_bits; // @[pearray.scala 156:36]
  assign PENetwork_36_io_to_pes_2_out_bits = PE_20_io_data_2_out_bits; // @[pearray.scala 156:36]
  assign PENetwork_36_io_to_pes_3_out_bits = PE_28_io_data_2_out_bits; // @[pearray.scala 156:36]
  assign PENetwork_36_io_to_pes_4_out_bits = PE_36_io_data_2_out_bits; // @[pearray.scala 156:36]
  assign PENetwork_36_io_to_pes_5_out_bits = PE_44_io_data_2_out_bits; // @[pearray.scala 156:36]
  assign PENetwork_36_io_to_pes_6_out_bits = PE_52_io_data_2_out_bits; // @[pearray.scala 156:36]
  assign PENetwork_36_io_to_pes_7_out_bits = PE_60_io_data_2_out_bits; // @[pearray.scala 156:36]
  assign PENetwork_36_io_to_pes_8_out_bits = PE_68_io_data_2_out_bits; // @[pearray.scala 156:36]
  assign PENetwork_36_io_to_pes_9_out_bits = PE_76_io_data_2_out_bits; // @[pearray.scala 156:36]
  assign PENetwork_36_io_to_pes_10_out_bits = PE_84_io_data_2_out_bits; // @[pearray.scala 156:36]
  assign PENetwork_36_io_to_pes_11_out_bits = PE_92_io_data_2_out_bits; // @[pearray.scala 156:36]
  assign PENetwork_36_io_to_pes_12_out_bits = PE_100_io_data_2_out_bits; // @[pearray.scala 156:36]
  assign PENetwork_36_io_to_pes_13_out_bits = PE_108_io_data_2_out_bits; // @[pearray.scala 156:36]
  assign PENetwork_36_io_to_pes_14_out_bits = PE_116_io_data_2_out_bits; // @[pearray.scala 156:36]
  assign PENetwork_36_io_to_mem_bits = MemController_36_io_rd_data_bits; // @[pearray.scala 239:29]
  assign PENetwork_37_io_to_pes_0_out_bits = PE_5_io_data_2_out_bits; // @[pearray.scala 156:36]
  assign PENetwork_37_io_to_pes_1_out_bits = PE_13_io_data_2_out_bits; // @[pearray.scala 156:36]
  assign PENetwork_37_io_to_pes_2_out_bits = PE_21_io_data_2_out_bits; // @[pearray.scala 156:36]
  assign PENetwork_37_io_to_pes_3_out_bits = PE_29_io_data_2_out_bits; // @[pearray.scala 156:36]
  assign PENetwork_37_io_to_pes_4_out_bits = PE_37_io_data_2_out_bits; // @[pearray.scala 156:36]
  assign PENetwork_37_io_to_pes_5_out_bits = PE_45_io_data_2_out_bits; // @[pearray.scala 156:36]
  assign PENetwork_37_io_to_pes_6_out_bits = PE_53_io_data_2_out_bits; // @[pearray.scala 156:36]
  assign PENetwork_37_io_to_pes_7_out_bits = PE_61_io_data_2_out_bits; // @[pearray.scala 156:36]
  assign PENetwork_37_io_to_pes_8_out_bits = PE_69_io_data_2_out_bits; // @[pearray.scala 156:36]
  assign PENetwork_37_io_to_pes_9_out_bits = PE_77_io_data_2_out_bits; // @[pearray.scala 156:36]
  assign PENetwork_37_io_to_pes_10_out_bits = PE_85_io_data_2_out_bits; // @[pearray.scala 156:36]
  assign PENetwork_37_io_to_pes_11_out_bits = PE_93_io_data_2_out_bits; // @[pearray.scala 156:36]
  assign PENetwork_37_io_to_pes_12_out_bits = PE_101_io_data_2_out_bits; // @[pearray.scala 156:36]
  assign PENetwork_37_io_to_pes_13_out_bits = PE_109_io_data_2_out_bits; // @[pearray.scala 156:36]
  assign PENetwork_37_io_to_pes_14_out_bits = PE_117_io_data_2_out_bits; // @[pearray.scala 156:36]
  assign PENetwork_37_io_to_mem_bits = MemController_37_io_rd_data_bits; // @[pearray.scala 239:29]
  assign PENetwork_38_io_to_pes_0_out_bits = PE_6_io_data_2_out_bits; // @[pearray.scala 156:36]
  assign PENetwork_38_io_to_pes_1_out_bits = PE_14_io_data_2_out_bits; // @[pearray.scala 156:36]
  assign PENetwork_38_io_to_pes_2_out_bits = PE_22_io_data_2_out_bits; // @[pearray.scala 156:36]
  assign PENetwork_38_io_to_pes_3_out_bits = PE_30_io_data_2_out_bits; // @[pearray.scala 156:36]
  assign PENetwork_38_io_to_pes_4_out_bits = PE_38_io_data_2_out_bits; // @[pearray.scala 156:36]
  assign PENetwork_38_io_to_pes_5_out_bits = PE_46_io_data_2_out_bits; // @[pearray.scala 156:36]
  assign PENetwork_38_io_to_pes_6_out_bits = PE_54_io_data_2_out_bits; // @[pearray.scala 156:36]
  assign PENetwork_38_io_to_pes_7_out_bits = PE_62_io_data_2_out_bits; // @[pearray.scala 156:36]
  assign PENetwork_38_io_to_pes_8_out_bits = PE_70_io_data_2_out_bits; // @[pearray.scala 156:36]
  assign PENetwork_38_io_to_pes_9_out_bits = PE_78_io_data_2_out_bits; // @[pearray.scala 156:36]
  assign PENetwork_38_io_to_pes_10_out_bits = PE_86_io_data_2_out_bits; // @[pearray.scala 156:36]
  assign PENetwork_38_io_to_pes_11_out_bits = PE_94_io_data_2_out_bits; // @[pearray.scala 156:36]
  assign PENetwork_38_io_to_pes_12_out_bits = PE_102_io_data_2_out_bits; // @[pearray.scala 156:36]
  assign PENetwork_38_io_to_pes_13_out_bits = PE_110_io_data_2_out_bits; // @[pearray.scala 156:36]
  assign PENetwork_38_io_to_pes_14_out_bits = PE_118_io_data_2_out_bits; // @[pearray.scala 156:36]
  assign PENetwork_38_io_to_mem_bits = MemController_38_io_rd_data_bits; // @[pearray.scala 239:29]
  assign PENetwork_39_io_to_pes_0_out_bits = PE_7_io_data_2_out_bits; // @[pearray.scala 156:36]
  assign PENetwork_39_io_to_pes_1_out_bits = PE_15_io_data_2_out_bits; // @[pearray.scala 156:36]
  assign PENetwork_39_io_to_pes_2_out_bits = PE_23_io_data_2_out_bits; // @[pearray.scala 156:36]
  assign PENetwork_39_io_to_pes_3_out_bits = PE_31_io_data_2_out_bits; // @[pearray.scala 156:36]
  assign PENetwork_39_io_to_pes_4_out_bits = PE_39_io_data_2_out_bits; // @[pearray.scala 156:36]
  assign PENetwork_39_io_to_pes_5_out_bits = PE_47_io_data_2_out_bits; // @[pearray.scala 156:36]
  assign PENetwork_39_io_to_pes_6_out_bits = PE_55_io_data_2_out_bits; // @[pearray.scala 156:36]
  assign PENetwork_39_io_to_pes_7_out_bits = PE_63_io_data_2_out_bits; // @[pearray.scala 156:36]
  assign PENetwork_39_io_to_pes_8_out_bits = PE_71_io_data_2_out_bits; // @[pearray.scala 156:36]
  assign PENetwork_39_io_to_pes_9_out_bits = PE_79_io_data_2_out_bits; // @[pearray.scala 156:36]
  assign PENetwork_39_io_to_pes_10_out_bits = PE_87_io_data_2_out_bits; // @[pearray.scala 156:36]
  assign PENetwork_39_io_to_pes_11_out_bits = PE_95_io_data_2_out_bits; // @[pearray.scala 156:36]
  assign PENetwork_39_io_to_pes_12_out_bits = PE_103_io_data_2_out_bits; // @[pearray.scala 156:36]
  assign PENetwork_39_io_to_pes_13_out_bits = PE_111_io_data_2_out_bits; // @[pearray.scala 156:36]
  assign PENetwork_39_io_to_pes_14_out_bits = PE_119_io_data_2_out_bits; // @[pearray.scala 156:36]
  assign PENetwork_39_io_to_mem_bits = MemController_39_io_rd_data_bits; // @[pearray.scala 239:29]
  assign MemController_clock = clock;
  assign MemController_reset = reset;
  assign MemController_io_rd_valid = io_out_valid; // @[pearray.scala 242:28]
  assign MemController_io_wr_valid = PENetwork_io_to_mem_valid; // @[pearray.scala 241:28]
  assign MemController_io_wr_data_valid = PENetwork_io_to_mem_valid; // @[pearray.scala 243:27]
  assign MemController_io_wr_data_bits = PENetwork_io_to_mem_bits; // @[pearray.scala 243:27]
  assign MemController_1_clock = clock;
  assign MemController_1_reset = reset;
  assign MemController_1_io_rd_valid = io_out_valid; // @[pearray.scala 242:28]
  assign MemController_1_io_wr_valid = PENetwork_1_io_to_mem_valid; // @[pearray.scala 241:28]
  assign MemController_1_io_wr_data_valid = PENetwork_1_io_to_mem_valid; // @[pearray.scala 243:27]
  assign MemController_1_io_wr_data_bits = PENetwork_1_io_to_mem_bits; // @[pearray.scala 243:27]
  assign MemController_2_clock = clock;
  assign MemController_2_reset = reset;
  assign MemController_2_io_rd_valid = io_out_valid; // @[pearray.scala 242:28]
  assign MemController_2_io_wr_valid = PENetwork_2_io_to_mem_valid; // @[pearray.scala 241:28]
  assign MemController_2_io_wr_data_valid = PENetwork_2_io_to_mem_valid; // @[pearray.scala 243:27]
  assign MemController_2_io_wr_data_bits = PENetwork_2_io_to_mem_bits; // @[pearray.scala 243:27]
  assign MemController_3_clock = clock;
  assign MemController_3_reset = reset;
  assign MemController_3_io_rd_valid = io_out_valid; // @[pearray.scala 242:28]
  assign MemController_3_io_wr_valid = PENetwork_3_io_to_mem_valid; // @[pearray.scala 241:28]
  assign MemController_3_io_wr_data_valid = PENetwork_3_io_to_mem_valid; // @[pearray.scala 243:27]
  assign MemController_3_io_wr_data_bits = PENetwork_3_io_to_mem_bits; // @[pearray.scala 243:27]
  assign MemController_4_clock = clock;
  assign MemController_4_reset = reset;
  assign MemController_4_io_rd_valid = io_out_valid; // @[pearray.scala 242:28]
  assign MemController_4_io_wr_valid = PENetwork_4_io_to_mem_valid; // @[pearray.scala 241:28]
  assign MemController_4_io_wr_data_valid = PENetwork_4_io_to_mem_valid; // @[pearray.scala 243:27]
  assign MemController_4_io_wr_data_bits = PENetwork_4_io_to_mem_bits; // @[pearray.scala 243:27]
  assign MemController_5_clock = clock;
  assign MemController_5_reset = reset;
  assign MemController_5_io_rd_valid = io_out_valid; // @[pearray.scala 242:28]
  assign MemController_5_io_wr_valid = PENetwork_5_io_to_mem_valid; // @[pearray.scala 241:28]
  assign MemController_5_io_wr_data_valid = PENetwork_5_io_to_mem_valid; // @[pearray.scala 243:27]
  assign MemController_5_io_wr_data_bits = PENetwork_5_io_to_mem_bits; // @[pearray.scala 243:27]
  assign MemController_6_clock = clock;
  assign MemController_6_reset = reset;
  assign MemController_6_io_rd_valid = io_out_valid; // @[pearray.scala 242:28]
  assign MemController_6_io_wr_valid = PENetwork_6_io_to_mem_valid; // @[pearray.scala 241:28]
  assign MemController_6_io_wr_data_valid = PENetwork_6_io_to_mem_valid; // @[pearray.scala 243:27]
  assign MemController_6_io_wr_data_bits = PENetwork_6_io_to_mem_bits; // @[pearray.scala 243:27]
  assign MemController_7_clock = clock;
  assign MemController_7_reset = reset;
  assign MemController_7_io_rd_valid = io_out_valid; // @[pearray.scala 242:28]
  assign MemController_7_io_wr_valid = PENetwork_7_io_to_mem_valid; // @[pearray.scala 241:28]
  assign MemController_7_io_wr_data_valid = PENetwork_7_io_to_mem_valid; // @[pearray.scala 243:27]
  assign MemController_7_io_wr_data_bits = PENetwork_7_io_to_mem_bits; // @[pearray.scala 243:27]
  assign MemController_8_clock = clock;
  assign MemController_8_reset = reset;
  assign MemController_8_io_rd_valid = io_out_valid; // @[pearray.scala 242:28]
  assign MemController_8_io_wr_valid = PENetwork_8_io_to_mem_valid; // @[pearray.scala 241:28]
  assign MemController_8_io_wr_data_valid = PENetwork_8_io_to_mem_valid; // @[pearray.scala 243:27]
  assign MemController_8_io_wr_data_bits = PENetwork_8_io_to_mem_bits; // @[pearray.scala 243:27]
  assign MemController_9_clock = clock;
  assign MemController_9_reset = reset;
  assign MemController_9_io_rd_valid = io_out_valid; // @[pearray.scala 242:28]
  assign MemController_9_io_wr_valid = PENetwork_9_io_to_mem_valid; // @[pearray.scala 241:28]
  assign MemController_9_io_wr_data_valid = PENetwork_9_io_to_mem_valid; // @[pearray.scala 243:27]
  assign MemController_9_io_wr_data_bits = PENetwork_9_io_to_mem_bits; // @[pearray.scala 243:27]
  assign MemController_10_clock = clock;
  assign MemController_10_reset = reset;
  assign MemController_10_io_rd_valid = io_out_valid; // @[pearray.scala 242:28]
  assign MemController_10_io_wr_valid = PENetwork_10_io_to_mem_valid; // @[pearray.scala 241:28]
  assign MemController_10_io_wr_data_valid = PENetwork_10_io_to_mem_valid; // @[pearray.scala 243:27]
  assign MemController_10_io_wr_data_bits = PENetwork_10_io_to_mem_bits; // @[pearray.scala 243:27]
  assign MemController_11_clock = clock;
  assign MemController_11_reset = reset;
  assign MemController_11_io_rd_valid = io_out_valid; // @[pearray.scala 242:28]
  assign MemController_11_io_wr_valid = PENetwork_11_io_to_mem_valid; // @[pearray.scala 241:28]
  assign MemController_11_io_wr_data_valid = PENetwork_11_io_to_mem_valid; // @[pearray.scala 243:27]
  assign MemController_11_io_wr_data_bits = PENetwork_11_io_to_mem_bits; // @[pearray.scala 243:27]
  assign MemController_12_clock = clock;
  assign MemController_12_reset = reset;
  assign MemController_12_io_rd_valid = io_out_valid; // @[pearray.scala 242:28]
  assign MemController_12_io_wr_valid = PENetwork_12_io_to_mem_valid; // @[pearray.scala 241:28]
  assign MemController_12_io_wr_data_valid = PENetwork_12_io_to_mem_valid; // @[pearray.scala 243:27]
  assign MemController_12_io_wr_data_bits = PENetwork_12_io_to_mem_bits; // @[pearray.scala 243:27]
  assign MemController_13_clock = clock;
  assign MemController_13_reset = reset;
  assign MemController_13_io_rd_valid = io_out_valid; // @[pearray.scala 242:28]
  assign MemController_13_io_wr_valid = PENetwork_13_io_to_mem_valid; // @[pearray.scala 241:28]
  assign MemController_13_io_wr_data_valid = PENetwork_13_io_to_mem_valid; // @[pearray.scala 243:27]
  assign MemController_13_io_wr_data_bits = PENetwork_13_io_to_mem_bits; // @[pearray.scala 243:27]
  assign MemController_14_clock = clock;
  assign MemController_14_reset = reset;
  assign MemController_14_io_rd_valid = io_out_valid; // @[pearray.scala 242:28]
  assign MemController_14_io_wr_valid = PENetwork_14_io_to_mem_valid; // @[pearray.scala 241:28]
  assign MemController_14_io_wr_data_valid = PENetwork_14_io_to_mem_valid; // @[pearray.scala 243:27]
  assign MemController_14_io_wr_data_bits = PENetwork_14_io_to_mem_bits; // @[pearray.scala 243:27]
  assign MemController_15_clock = clock;
  assign MemController_15_reset = reset;
  assign MemController_15_io_rd_valid = io_out_valid; // @[pearray.scala 242:28]
  assign MemController_15_io_wr_valid = PENetwork_15_io_to_mem_valid; // @[pearray.scala 241:28]
  assign MemController_15_io_wr_data_valid = PENetwork_15_io_to_mem_valid; // @[pearray.scala 243:27]
  assign MemController_15_io_wr_data_bits = PENetwork_15_io_to_mem_bits; // @[pearray.scala 243:27]
  assign MemController_16_clock = clock;
  assign MemController_16_reset = reset;
  assign MemController_16_io_rd_valid = _T_1585_2; // @[pearray.scala 236:30]
  assign MemController_16_io_wr_valid = io_data_1_in_0_valid; // @[pearray.scala 237:28]
  assign MemController_16_io_wr_data_valid = io_data_1_in_0_bits_valid; // @[pearray.scala 238:27]
  assign MemController_16_io_wr_data_bits = io_data_1_in_0_bits_bits; // @[pearray.scala 238:27]
  assign MemController_17_clock = clock;
  assign MemController_17_reset = reset;
  assign MemController_17_io_rd_valid = _T_1594_2; // @[pearray.scala 236:30]
  assign MemController_17_io_wr_valid = io_data_1_in_1_valid; // @[pearray.scala 237:28]
  assign MemController_17_io_wr_data_valid = io_data_1_in_1_bits_valid; // @[pearray.scala 238:27]
  assign MemController_17_io_wr_data_bits = io_data_1_in_1_bits_bits; // @[pearray.scala 238:27]
  assign MemController_18_clock = clock;
  assign MemController_18_reset = reset;
  assign MemController_18_io_rd_valid = _T_1603_2; // @[pearray.scala 236:30]
  assign MemController_18_io_wr_valid = io_data_1_in_2_valid; // @[pearray.scala 237:28]
  assign MemController_18_io_wr_data_valid = io_data_1_in_2_bits_valid; // @[pearray.scala 238:27]
  assign MemController_18_io_wr_data_bits = io_data_1_in_2_bits_bits; // @[pearray.scala 238:27]
  assign MemController_19_clock = clock;
  assign MemController_19_reset = reset;
  assign MemController_19_io_rd_valid = _T_1612_2; // @[pearray.scala 236:30]
  assign MemController_19_io_wr_valid = io_data_1_in_3_valid; // @[pearray.scala 237:28]
  assign MemController_19_io_wr_data_valid = io_data_1_in_3_bits_valid; // @[pearray.scala 238:27]
  assign MemController_19_io_wr_data_bits = io_data_1_in_3_bits_bits; // @[pearray.scala 238:27]
  assign MemController_20_clock = clock;
  assign MemController_20_reset = reset;
  assign MemController_20_io_rd_valid = _T_1621_2; // @[pearray.scala 236:30]
  assign MemController_20_io_wr_valid = io_data_1_in_4_valid; // @[pearray.scala 237:28]
  assign MemController_20_io_wr_data_valid = io_data_1_in_4_bits_valid; // @[pearray.scala 238:27]
  assign MemController_20_io_wr_data_bits = io_data_1_in_4_bits_bits; // @[pearray.scala 238:27]
  assign MemController_21_clock = clock;
  assign MemController_21_reset = reset;
  assign MemController_21_io_rd_valid = _T_1630_2; // @[pearray.scala 236:30]
  assign MemController_21_io_wr_valid = io_data_1_in_5_valid; // @[pearray.scala 237:28]
  assign MemController_21_io_wr_data_valid = io_data_1_in_5_bits_valid; // @[pearray.scala 238:27]
  assign MemController_21_io_wr_data_bits = io_data_1_in_5_bits_bits; // @[pearray.scala 238:27]
  assign MemController_22_clock = clock;
  assign MemController_22_reset = reset;
  assign MemController_22_io_rd_valid = _T_1639_2; // @[pearray.scala 236:30]
  assign MemController_22_io_wr_valid = io_data_1_in_6_valid; // @[pearray.scala 237:28]
  assign MemController_22_io_wr_data_valid = io_data_1_in_6_bits_valid; // @[pearray.scala 238:27]
  assign MemController_22_io_wr_data_bits = io_data_1_in_6_bits_bits; // @[pearray.scala 238:27]
  assign MemController_23_clock = clock;
  assign MemController_23_reset = reset;
  assign MemController_23_io_rd_valid = _T_1648_2; // @[pearray.scala 236:30]
  assign MemController_23_io_wr_valid = io_data_1_in_7_valid; // @[pearray.scala 237:28]
  assign MemController_23_io_wr_data_valid = io_data_1_in_7_bits_valid; // @[pearray.scala 238:27]
  assign MemController_23_io_wr_data_bits = io_data_1_in_7_bits_bits; // @[pearray.scala 238:27]
  assign MemController_24_clock = clock;
  assign MemController_24_reset = reset;
  assign MemController_24_io_rd_valid = _T_1657_2; // @[pearray.scala 236:30]
  assign MemController_24_io_wr_valid = io_data_1_in_8_valid; // @[pearray.scala 237:28]
  assign MemController_24_io_wr_data_valid = io_data_1_in_8_bits_valid; // @[pearray.scala 238:27]
  assign MemController_24_io_wr_data_bits = io_data_1_in_8_bits_bits; // @[pearray.scala 238:27]
  assign MemController_25_clock = clock;
  assign MemController_25_reset = reset;
  assign MemController_25_io_rd_valid = _T_1666_2; // @[pearray.scala 236:30]
  assign MemController_25_io_wr_valid = io_data_1_in_9_valid; // @[pearray.scala 237:28]
  assign MemController_25_io_wr_data_valid = io_data_1_in_9_bits_valid; // @[pearray.scala 238:27]
  assign MemController_25_io_wr_data_bits = io_data_1_in_9_bits_bits; // @[pearray.scala 238:27]
  assign MemController_26_clock = clock;
  assign MemController_26_reset = reset;
  assign MemController_26_io_rd_valid = _T_1675_2; // @[pearray.scala 236:30]
  assign MemController_26_io_wr_valid = io_data_1_in_10_valid; // @[pearray.scala 237:28]
  assign MemController_26_io_wr_data_valid = io_data_1_in_10_bits_valid; // @[pearray.scala 238:27]
  assign MemController_26_io_wr_data_bits = io_data_1_in_10_bits_bits; // @[pearray.scala 238:27]
  assign MemController_27_clock = clock;
  assign MemController_27_reset = reset;
  assign MemController_27_io_rd_valid = _T_1684_2; // @[pearray.scala 236:30]
  assign MemController_27_io_wr_valid = io_data_1_in_11_valid; // @[pearray.scala 237:28]
  assign MemController_27_io_wr_data_valid = io_data_1_in_11_bits_valid; // @[pearray.scala 238:27]
  assign MemController_27_io_wr_data_bits = io_data_1_in_11_bits_bits; // @[pearray.scala 238:27]
  assign MemController_28_clock = clock;
  assign MemController_28_reset = reset;
  assign MemController_28_io_rd_valid = _T_1693_2; // @[pearray.scala 236:30]
  assign MemController_28_io_wr_valid = io_data_1_in_12_valid; // @[pearray.scala 237:28]
  assign MemController_28_io_wr_data_valid = io_data_1_in_12_bits_valid; // @[pearray.scala 238:27]
  assign MemController_28_io_wr_data_bits = io_data_1_in_12_bits_bits; // @[pearray.scala 238:27]
  assign MemController_29_clock = clock;
  assign MemController_29_reset = reset;
  assign MemController_29_io_rd_valid = _T_1702_2; // @[pearray.scala 236:30]
  assign MemController_29_io_wr_valid = io_data_1_in_13_valid; // @[pearray.scala 237:28]
  assign MemController_29_io_wr_data_valid = io_data_1_in_13_bits_valid; // @[pearray.scala 238:27]
  assign MemController_29_io_wr_data_bits = io_data_1_in_13_bits_bits; // @[pearray.scala 238:27]
  assign MemController_30_clock = clock;
  assign MemController_30_reset = reset;
  assign MemController_30_io_rd_valid = _T_1711_2; // @[pearray.scala 236:30]
  assign MemController_30_io_wr_valid = io_data_1_in_14_valid; // @[pearray.scala 237:28]
  assign MemController_30_io_wr_data_valid = io_data_1_in_14_bits_valid; // @[pearray.scala 238:27]
  assign MemController_30_io_wr_data_bits = io_data_1_in_14_bits_bits; // @[pearray.scala 238:27]
  assign MemController_31_clock = clock;
  assign MemController_31_reset = reset;
  assign MemController_31_io_rd_valid = _T_1720_2; // @[pearray.scala 236:30]
  assign MemController_31_io_wr_valid = io_data_1_in_15_valid; // @[pearray.scala 237:28]
  assign MemController_31_io_wr_data_valid = io_data_1_in_15_bits_valid; // @[pearray.scala 238:27]
  assign MemController_31_io_wr_data_bits = io_data_1_in_15_bits_bits; // @[pearray.scala 238:27]
  assign MemController_32_clock = clock;
  assign MemController_32_reset = reset;
  assign MemController_32_io_rd_valid = io_exec_valid; // @[pearray.scala 229:32]
  assign MemController_32_io_wr_valid = io_data_2_in_0_valid; // @[pearray.scala 237:28]
  assign MemController_32_io_wr_data_valid = io_data_2_in_0_bits_valid; // @[pearray.scala 238:27]
  assign MemController_32_io_wr_data_bits = io_data_2_in_0_bits_bits; // @[pearray.scala 238:27]
  assign MemController_33_clock = clock;
  assign MemController_33_reset = reset;
  assign MemController_33_io_rd_valid = _T_1722_0; // @[pearray.scala 227:32]
  assign MemController_33_io_wr_valid = io_data_2_in_1_valid; // @[pearray.scala 237:28]
  assign MemController_33_io_wr_data_valid = io_data_2_in_1_bits_valid; // @[pearray.scala 238:27]
  assign MemController_33_io_wr_data_bits = io_data_2_in_1_bits_bits; // @[pearray.scala 238:27]
  assign MemController_34_clock = clock;
  assign MemController_34_reset = reset;
  assign MemController_34_io_rd_valid = _T_1722_1; // @[pearray.scala 227:32]
  assign MemController_34_io_wr_valid = io_data_2_in_2_valid; // @[pearray.scala 237:28]
  assign MemController_34_io_wr_data_valid = io_data_2_in_2_bits_valid; // @[pearray.scala 238:27]
  assign MemController_34_io_wr_data_bits = io_data_2_in_2_bits_bits; // @[pearray.scala 238:27]
  assign MemController_35_clock = clock;
  assign MemController_35_reset = reset;
  assign MemController_35_io_rd_valid = _T_1722_2; // @[pearray.scala 227:32]
  assign MemController_35_io_wr_valid = io_data_2_in_3_valid; // @[pearray.scala 237:28]
  assign MemController_35_io_wr_data_valid = io_data_2_in_3_bits_valid; // @[pearray.scala 238:27]
  assign MemController_35_io_wr_data_bits = io_data_2_in_3_bits_bits; // @[pearray.scala 238:27]
  assign MemController_36_clock = clock;
  assign MemController_36_reset = reset;
  assign MemController_36_io_rd_valid = _T_1722_3; // @[pearray.scala 227:32]
  assign MemController_36_io_wr_valid = io_data_2_in_4_valid; // @[pearray.scala 237:28]
  assign MemController_36_io_wr_data_valid = io_data_2_in_4_bits_valid; // @[pearray.scala 238:27]
  assign MemController_36_io_wr_data_bits = io_data_2_in_4_bits_bits; // @[pearray.scala 238:27]
  assign MemController_37_clock = clock;
  assign MemController_37_reset = reset;
  assign MemController_37_io_rd_valid = _T_1722_4; // @[pearray.scala 227:32]
  assign MemController_37_io_wr_valid = io_data_2_in_5_valid; // @[pearray.scala 237:28]
  assign MemController_37_io_wr_data_valid = io_data_2_in_5_bits_valid; // @[pearray.scala 238:27]
  assign MemController_37_io_wr_data_bits = io_data_2_in_5_bits_bits; // @[pearray.scala 238:27]
  assign MemController_38_clock = clock;
  assign MemController_38_reset = reset;
  assign MemController_38_io_rd_valid = _T_1722_5; // @[pearray.scala 227:32]
  assign MemController_38_io_wr_valid = io_data_2_in_6_valid; // @[pearray.scala 237:28]
  assign MemController_38_io_wr_data_valid = io_data_2_in_6_bits_valid; // @[pearray.scala 238:27]
  assign MemController_38_io_wr_data_bits = io_data_2_in_6_bits_bits; // @[pearray.scala 238:27]
  assign MemController_39_clock = clock;
  assign MemController_39_reset = reset;
  assign MemController_39_io_rd_valid = _T_1722_6; // @[pearray.scala 227:32]
  assign MemController_39_io_wr_valid = io_data_2_in_7_valid; // @[pearray.scala 237:28]
  assign MemController_39_io_wr_data_valid = io_data_2_in_7_bits_valid; // @[pearray.scala 238:27]
  assign MemController_39_io_wr_data_bits = io_data_2_in_7_bits_bits; // @[pearray.scala 238:27]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _T_16_0 = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  _T_16_1 = _RAND_1[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  _T_16_2 = _RAND_2[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  _T_16_3 = _RAND_3[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  _T_28_0 = _RAND_4[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{`RANDOM}};
  _T_28_1 = _RAND_5[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {1{`RANDOM}};
  _T_28_2 = _RAND_6[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7 = {1{`RANDOM}};
  _T_28_3 = _RAND_7[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8 = {1{`RANDOM}};
  _T_40_0 = _RAND_8[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9 = {1{`RANDOM}};
  _T_40_1 = _RAND_9[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10 = {1{`RANDOM}};
  _T_40_2 = _RAND_10[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11 = {1{`RANDOM}};
  _T_40_3 = _RAND_11[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_12 = {1{`RANDOM}};
  _T_52_0 = _RAND_12[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_13 = {1{`RANDOM}};
  _T_52_1 = _RAND_13[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_14 = {1{`RANDOM}};
  _T_52_2 = _RAND_14[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_15 = {1{`RANDOM}};
  _T_52_3 = _RAND_15[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_16 = {1{`RANDOM}};
  _T_64_0 = _RAND_16[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_17 = {1{`RANDOM}};
  _T_64_1 = _RAND_17[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_18 = {1{`RANDOM}};
  _T_64_2 = _RAND_18[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_19 = {1{`RANDOM}};
  _T_64_3 = _RAND_19[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_20 = {1{`RANDOM}};
  _T_76_0 = _RAND_20[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_21 = {1{`RANDOM}};
  _T_76_1 = _RAND_21[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_22 = {1{`RANDOM}};
  _T_76_2 = _RAND_22[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_23 = {1{`RANDOM}};
  _T_76_3 = _RAND_23[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_24 = {1{`RANDOM}};
  _T_88_0 = _RAND_24[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_25 = {1{`RANDOM}};
  _T_88_1 = _RAND_25[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_26 = {1{`RANDOM}};
  _T_88_2 = _RAND_26[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_27 = {1{`RANDOM}};
  _T_88_3 = _RAND_27[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_28 = {1{`RANDOM}};
  _T_100_0 = _RAND_28[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_29 = {1{`RANDOM}};
  _T_100_1 = _RAND_29[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_30 = {1{`RANDOM}};
  _T_100_2 = _RAND_30[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_31 = {1{`RANDOM}};
  _T_100_3 = _RAND_31[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_32 = {1{`RANDOM}};
  _T_114_0 = _RAND_32[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_33 = {1{`RANDOM}};
  _T_114_1 = _RAND_33[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_34 = {1{`RANDOM}};
  _T_114_2 = _RAND_34[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_35 = {1{`RANDOM}};
  _T_114_3 = _RAND_35[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_36 = {1{`RANDOM}};
  _T_126_0 = _RAND_36[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_37 = {1{`RANDOM}};
  _T_126_1 = _RAND_37[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_38 = {1{`RANDOM}};
  _T_126_2 = _RAND_38[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_39 = {1{`RANDOM}};
  _T_126_3 = _RAND_39[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_40 = {1{`RANDOM}};
  _T_138_0 = _RAND_40[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_41 = {1{`RANDOM}};
  _T_138_1 = _RAND_41[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_42 = {1{`RANDOM}};
  _T_138_2 = _RAND_42[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_43 = {1{`RANDOM}};
  _T_138_3 = _RAND_43[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_44 = {1{`RANDOM}};
  _T_150_0 = _RAND_44[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_45 = {1{`RANDOM}};
  _T_150_1 = _RAND_45[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_46 = {1{`RANDOM}};
  _T_150_2 = _RAND_46[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_47 = {1{`RANDOM}};
  _T_150_3 = _RAND_47[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_48 = {1{`RANDOM}};
  _T_162_0 = _RAND_48[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_49 = {1{`RANDOM}};
  _T_162_1 = _RAND_49[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_50 = {1{`RANDOM}};
  _T_162_2 = _RAND_50[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_51 = {1{`RANDOM}};
  _T_162_3 = _RAND_51[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_52 = {1{`RANDOM}};
  _T_174_0 = _RAND_52[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_53 = {1{`RANDOM}};
  _T_174_1 = _RAND_53[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_54 = {1{`RANDOM}};
  _T_174_2 = _RAND_54[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_55 = {1{`RANDOM}};
  _T_174_3 = _RAND_55[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_56 = {1{`RANDOM}};
  _T_186_0 = _RAND_56[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_57 = {1{`RANDOM}};
  _T_186_1 = _RAND_57[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_58 = {1{`RANDOM}};
  _T_186_2 = _RAND_58[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_59 = {1{`RANDOM}};
  _T_186_3 = _RAND_59[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_60 = {1{`RANDOM}};
  _T_198_0 = _RAND_60[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_61 = {1{`RANDOM}};
  _T_198_1 = _RAND_61[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_62 = {1{`RANDOM}};
  _T_198_2 = _RAND_62[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_63 = {1{`RANDOM}};
  _T_198_3 = _RAND_63[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_64 = {1{`RANDOM}};
  _T_212_0 = _RAND_64[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_65 = {1{`RANDOM}};
  _T_212_1 = _RAND_65[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_66 = {1{`RANDOM}};
  _T_212_2 = _RAND_66[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_67 = {1{`RANDOM}};
  _T_212_3 = _RAND_67[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_68 = {1{`RANDOM}};
  _T_224_0 = _RAND_68[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_69 = {1{`RANDOM}};
  _T_224_1 = _RAND_69[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_70 = {1{`RANDOM}};
  _T_224_2 = _RAND_70[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_71 = {1{`RANDOM}};
  _T_224_3 = _RAND_71[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_72 = {1{`RANDOM}};
  _T_236_0 = _RAND_72[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_73 = {1{`RANDOM}};
  _T_236_1 = _RAND_73[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_74 = {1{`RANDOM}};
  _T_236_2 = _RAND_74[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_75 = {1{`RANDOM}};
  _T_236_3 = _RAND_75[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_76 = {1{`RANDOM}};
  _T_248_0 = _RAND_76[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_77 = {1{`RANDOM}};
  _T_248_1 = _RAND_77[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_78 = {1{`RANDOM}};
  _T_248_2 = _RAND_78[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_79 = {1{`RANDOM}};
  _T_248_3 = _RAND_79[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_80 = {1{`RANDOM}};
  _T_260_0 = _RAND_80[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_81 = {1{`RANDOM}};
  _T_260_1 = _RAND_81[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_82 = {1{`RANDOM}};
  _T_260_2 = _RAND_82[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_83 = {1{`RANDOM}};
  _T_260_3 = _RAND_83[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_84 = {1{`RANDOM}};
  _T_272_0 = _RAND_84[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_85 = {1{`RANDOM}};
  _T_272_1 = _RAND_85[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_86 = {1{`RANDOM}};
  _T_272_2 = _RAND_86[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_87 = {1{`RANDOM}};
  _T_272_3 = _RAND_87[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_88 = {1{`RANDOM}};
  _T_284_0 = _RAND_88[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_89 = {1{`RANDOM}};
  _T_284_1 = _RAND_89[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_90 = {1{`RANDOM}};
  _T_284_2 = _RAND_90[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_91 = {1{`RANDOM}};
  _T_284_3 = _RAND_91[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_92 = {1{`RANDOM}};
  _T_296_0 = _RAND_92[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_93 = {1{`RANDOM}};
  _T_296_1 = _RAND_93[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_94 = {1{`RANDOM}};
  _T_296_2 = _RAND_94[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_95 = {1{`RANDOM}};
  _T_296_3 = _RAND_95[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_96 = {1{`RANDOM}};
  _T_310_0 = _RAND_96[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_97 = {1{`RANDOM}};
  _T_310_1 = _RAND_97[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_98 = {1{`RANDOM}};
  _T_310_2 = _RAND_98[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_99 = {1{`RANDOM}};
  _T_310_3 = _RAND_99[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_100 = {1{`RANDOM}};
  _T_322_0 = _RAND_100[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_101 = {1{`RANDOM}};
  _T_322_1 = _RAND_101[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_102 = {1{`RANDOM}};
  _T_322_2 = _RAND_102[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_103 = {1{`RANDOM}};
  _T_322_3 = _RAND_103[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_104 = {1{`RANDOM}};
  _T_334_0 = _RAND_104[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_105 = {1{`RANDOM}};
  _T_334_1 = _RAND_105[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_106 = {1{`RANDOM}};
  _T_334_2 = _RAND_106[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_107 = {1{`RANDOM}};
  _T_334_3 = _RAND_107[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_108 = {1{`RANDOM}};
  _T_346_0 = _RAND_108[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_109 = {1{`RANDOM}};
  _T_346_1 = _RAND_109[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_110 = {1{`RANDOM}};
  _T_346_2 = _RAND_110[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_111 = {1{`RANDOM}};
  _T_346_3 = _RAND_111[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_112 = {1{`RANDOM}};
  _T_358_0 = _RAND_112[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_113 = {1{`RANDOM}};
  _T_358_1 = _RAND_113[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_114 = {1{`RANDOM}};
  _T_358_2 = _RAND_114[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_115 = {1{`RANDOM}};
  _T_358_3 = _RAND_115[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_116 = {1{`RANDOM}};
  _T_370_0 = _RAND_116[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_117 = {1{`RANDOM}};
  _T_370_1 = _RAND_117[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_118 = {1{`RANDOM}};
  _T_370_2 = _RAND_118[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_119 = {1{`RANDOM}};
  _T_370_3 = _RAND_119[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_120 = {1{`RANDOM}};
  _T_382_0 = _RAND_120[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_121 = {1{`RANDOM}};
  _T_382_1 = _RAND_121[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_122 = {1{`RANDOM}};
  _T_382_2 = _RAND_122[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_123 = {1{`RANDOM}};
  _T_382_3 = _RAND_123[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_124 = {1{`RANDOM}};
  _T_394_0 = _RAND_124[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_125 = {1{`RANDOM}};
  _T_394_1 = _RAND_125[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_126 = {1{`RANDOM}};
  _T_394_2 = _RAND_126[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_127 = {1{`RANDOM}};
  _T_394_3 = _RAND_127[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_128 = {1{`RANDOM}};
  _T_408_0 = _RAND_128[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_129 = {1{`RANDOM}};
  _T_408_1 = _RAND_129[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_130 = {1{`RANDOM}};
  _T_408_2 = _RAND_130[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_131 = {1{`RANDOM}};
  _T_408_3 = _RAND_131[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_132 = {1{`RANDOM}};
  _T_420_0 = _RAND_132[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_133 = {1{`RANDOM}};
  _T_420_1 = _RAND_133[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_134 = {1{`RANDOM}};
  _T_420_2 = _RAND_134[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_135 = {1{`RANDOM}};
  _T_420_3 = _RAND_135[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_136 = {1{`RANDOM}};
  _T_432_0 = _RAND_136[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_137 = {1{`RANDOM}};
  _T_432_1 = _RAND_137[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_138 = {1{`RANDOM}};
  _T_432_2 = _RAND_138[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_139 = {1{`RANDOM}};
  _T_432_3 = _RAND_139[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_140 = {1{`RANDOM}};
  _T_444_0 = _RAND_140[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_141 = {1{`RANDOM}};
  _T_444_1 = _RAND_141[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_142 = {1{`RANDOM}};
  _T_444_2 = _RAND_142[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_143 = {1{`RANDOM}};
  _T_444_3 = _RAND_143[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_144 = {1{`RANDOM}};
  _T_456_0 = _RAND_144[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_145 = {1{`RANDOM}};
  _T_456_1 = _RAND_145[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_146 = {1{`RANDOM}};
  _T_456_2 = _RAND_146[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_147 = {1{`RANDOM}};
  _T_456_3 = _RAND_147[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_148 = {1{`RANDOM}};
  _T_468_0 = _RAND_148[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_149 = {1{`RANDOM}};
  _T_468_1 = _RAND_149[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_150 = {1{`RANDOM}};
  _T_468_2 = _RAND_150[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_151 = {1{`RANDOM}};
  _T_468_3 = _RAND_151[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_152 = {1{`RANDOM}};
  _T_480_0 = _RAND_152[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_153 = {1{`RANDOM}};
  _T_480_1 = _RAND_153[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_154 = {1{`RANDOM}};
  _T_480_2 = _RAND_154[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_155 = {1{`RANDOM}};
  _T_480_3 = _RAND_155[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_156 = {1{`RANDOM}};
  _T_492_0 = _RAND_156[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_157 = {1{`RANDOM}};
  _T_492_1 = _RAND_157[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_158 = {1{`RANDOM}};
  _T_492_2 = _RAND_158[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_159 = {1{`RANDOM}};
  _T_492_3 = _RAND_159[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_160 = {1{`RANDOM}};
  _T_506_0 = _RAND_160[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_161 = {1{`RANDOM}};
  _T_506_1 = _RAND_161[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_162 = {1{`RANDOM}};
  _T_506_2 = _RAND_162[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_163 = {1{`RANDOM}};
  _T_506_3 = _RAND_163[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_164 = {1{`RANDOM}};
  _T_518_0 = _RAND_164[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_165 = {1{`RANDOM}};
  _T_518_1 = _RAND_165[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_166 = {1{`RANDOM}};
  _T_518_2 = _RAND_166[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_167 = {1{`RANDOM}};
  _T_518_3 = _RAND_167[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_168 = {1{`RANDOM}};
  _T_530_0 = _RAND_168[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_169 = {1{`RANDOM}};
  _T_530_1 = _RAND_169[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_170 = {1{`RANDOM}};
  _T_530_2 = _RAND_170[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_171 = {1{`RANDOM}};
  _T_530_3 = _RAND_171[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_172 = {1{`RANDOM}};
  _T_542_0 = _RAND_172[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_173 = {1{`RANDOM}};
  _T_542_1 = _RAND_173[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_174 = {1{`RANDOM}};
  _T_542_2 = _RAND_174[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_175 = {1{`RANDOM}};
  _T_542_3 = _RAND_175[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_176 = {1{`RANDOM}};
  _T_554_0 = _RAND_176[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_177 = {1{`RANDOM}};
  _T_554_1 = _RAND_177[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_178 = {1{`RANDOM}};
  _T_554_2 = _RAND_178[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_179 = {1{`RANDOM}};
  _T_554_3 = _RAND_179[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_180 = {1{`RANDOM}};
  _T_566_0 = _RAND_180[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_181 = {1{`RANDOM}};
  _T_566_1 = _RAND_181[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_182 = {1{`RANDOM}};
  _T_566_2 = _RAND_182[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_183 = {1{`RANDOM}};
  _T_566_3 = _RAND_183[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_184 = {1{`RANDOM}};
  _T_578_0 = _RAND_184[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_185 = {1{`RANDOM}};
  _T_578_1 = _RAND_185[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_186 = {1{`RANDOM}};
  _T_578_2 = _RAND_186[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_187 = {1{`RANDOM}};
  _T_578_3 = _RAND_187[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_188 = {1{`RANDOM}};
  _T_590_0 = _RAND_188[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_189 = {1{`RANDOM}};
  _T_590_1 = _RAND_189[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_190 = {1{`RANDOM}};
  _T_590_2 = _RAND_190[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_191 = {1{`RANDOM}};
  _T_590_3 = _RAND_191[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_192 = {1{`RANDOM}};
  _T_604_0 = _RAND_192[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_193 = {1{`RANDOM}};
  _T_604_1 = _RAND_193[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_194 = {1{`RANDOM}};
  _T_604_2 = _RAND_194[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_195 = {1{`RANDOM}};
  _T_604_3 = _RAND_195[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_196 = {1{`RANDOM}};
  _T_616_0 = _RAND_196[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_197 = {1{`RANDOM}};
  _T_616_1 = _RAND_197[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_198 = {1{`RANDOM}};
  _T_616_2 = _RAND_198[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_199 = {1{`RANDOM}};
  _T_616_3 = _RAND_199[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_200 = {1{`RANDOM}};
  _T_628_0 = _RAND_200[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_201 = {1{`RANDOM}};
  _T_628_1 = _RAND_201[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_202 = {1{`RANDOM}};
  _T_628_2 = _RAND_202[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_203 = {1{`RANDOM}};
  _T_628_3 = _RAND_203[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_204 = {1{`RANDOM}};
  _T_640_0 = _RAND_204[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_205 = {1{`RANDOM}};
  _T_640_1 = _RAND_205[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_206 = {1{`RANDOM}};
  _T_640_2 = _RAND_206[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_207 = {1{`RANDOM}};
  _T_640_3 = _RAND_207[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_208 = {1{`RANDOM}};
  _T_652_0 = _RAND_208[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_209 = {1{`RANDOM}};
  _T_652_1 = _RAND_209[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_210 = {1{`RANDOM}};
  _T_652_2 = _RAND_210[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_211 = {1{`RANDOM}};
  _T_652_3 = _RAND_211[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_212 = {1{`RANDOM}};
  _T_664_0 = _RAND_212[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_213 = {1{`RANDOM}};
  _T_664_1 = _RAND_213[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_214 = {1{`RANDOM}};
  _T_664_2 = _RAND_214[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_215 = {1{`RANDOM}};
  _T_664_3 = _RAND_215[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_216 = {1{`RANDOM}};
  _T_676_0 = _RAND_216[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_217 = {1{`RANDOM}};
  _T_676_1 = _RAND_217[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_218 = {1{`RANDOM}};
  _T_676_2 = _RAND_218[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_219 = {1{`RANDOM}};
  _T_676_3 = _RAND_219[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_220 = {1{`RANDOM}};
  _T_688_0 = _RAND_220[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_221 = {1{`RANDOM}};
  _T_688_1 = _RAND_221[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_222 = {1{`RANDOM}};
  _T_688_2 = _RAND_222[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_223 = {1{`RANDOM}};
  _T_688_3 = _RAND_223[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_224 = {1{`RANDOM}};
  _T_702_0 = _RAND_224[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_225 = {1{`RANDOM}};
  _T_702_1 = _RAND_225[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_226 = {1{`RANDOM}};
  _T_702_2 = _RAND_226[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_227 = {1{`RANDOM}};
  _T_702_3 = _RAND_227[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_228 = {1{`RANDOM}};
  _T_714_0 = _RAND_228[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_229 = {1{`RANDOM}};
  _T_714_1 = _RAND_229[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_230 = {1{`RANDOM}};
  _T_714_2 = _RAND_230[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_231 = {1{`RANDOM}};
  _T_714_3 = _RAND_231[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_232 = {1{`RANDOM}};
  _T_726_0 = _RAND_232[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_233 = {1{`RANDOM}};
  _T_726_1 = _RAND_233[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_234 = {1{`RANDOM}};
  _T_726_2 = _RAND_234[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_235 = {1{`RANDOM}};
  _T_726_3 = _RAND_235[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_236 = {1{`RANDOM}};
  _T_738_0 = _RAND_236[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_237 = {1{`RANDOM}};
  _T_738_1 = _RAND_237[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_238 = {1{`RANDOM}};
  _T_738_2 = _RAND_238[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_239 = {1{`RANDOM}};
  _T_738_3 = _RAND_239[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_240 = {1{`RANDOM}};
  _T_750_0 = _RAND_240[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_241 = {1{`RANDOM}};
  _T_750_1 = _RAND_241[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_242 = {1{`RANDOM}};
  _T_750_2 = _RAND_242[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_243 = {1{`RANDOM}};
  _T_750_3 = _RAND_243[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_244 = {1{`RANDOM}};
  _T_762_0 = _RAND_244[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_245 = {1{`RANDOM}};
  _T_762_1 = _RAND_245[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_246 = {1{`RANDOM}};
  _T_762_2 = _RAND_246[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_247 = {1{`RANDOM}};
  _T_762_3 = _RAND_247[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_248 = {1{`RANDOM}};
  _T_774_0 = _RAND_248[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_249 = {1{`RANDOM}};
  _T_774_1 = _RAND_249[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_250 = {1{`RANDOM}};
  _T_774_2 = _RAND_250[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_251 = {1{`RANDOM}};
  _T_774_3 = _RAND_251[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_252 = {1{`RANDOM}};
  _T_786_0 = _RAND_252[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_253 = {1{`RANDOM}};
  _T_786_1 = _RAND_253[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_254 = {1{`RANDOM}};
  _T_786_2 = _RAND_254[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_255 = {1{`RANDOM}};
  _T_786_3 = _RAND_255[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_256 = {1{`RANDOM}};
  _T_800_0 = _RAND_256[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_257 = {1{`RANDOM}};
  _T_800_1 = _RAND_257[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_258 = {1{`RANDOM}};
  _T_800_2 = _RAND_258[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_259 = {1{`RANDOM}};
  _T_800_3 = _RAND_259[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_260 = {1{`RANDOM}};
  _T_812_0 = _RAND_260[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_261 = {1{`RANDOM}};
  _T_812_1 = _RAND_261[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_262 = {1{`RANDOM}};
  _T_812_2 = _RAND_262[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_263 = {1{`RANDOM}};
  _T_812_3 = _RAND_263[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_264 = {1{`RANDOM}};
  _T_824_0 = _RAND_264[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_265 = {1{`RANDOM}};
  _T_824_1 = _RAND_265[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_266 = {1{`RANDOM}};
  _T_824_2 = _RAND_266[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_267 = {1{`RANDOM}};
  _T_824_3 = _RAND_267[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_268 = {1{`RANDOM}};
  _T_836_0 = _RAND_268[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_269 = {1{`RANDOM}};
  _T_836_1 = _RAND_269[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_270 = {1{`RANDOM}};
  _T_836_2 = _RAND_270[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_271 = {1{`RANDOM}};
  _T_836_3 = _RAND_271[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_272 = {1{`RANDOM}};
  _T_848_0 = _RAND_272[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_273 = {1{`RANDOM}};
  _T_848_1 = _RAND_273[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_274 = {1{`RANDOM}};
  _T_848_2 = _RAND_274[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_275 = {1{`RANDOM}};
  _T_848_3 = _RAND_275[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_276 = {1{`RANDOM}};
  _T_860_0 = _RAND_276[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_277 = {1{`RANDOM}};
  _T_860_1 = _RAND_277[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_278 = {1{`RANDOM}};
  _T_860_2 = _RAND_278[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_279 = {1{`RANDOM}};
  _T_860_3 = _RAND_279[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_280 = {1{`RANDOM}};
  _T_872_0 = _RAND_280[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_281 = {1{`RANDOM}};
  _T_872_1 = _RAND_281[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_282 = {1{`RANDOM}};
  _T_872_2 = _RAND_282[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_283 = {1{`RANDOM}};
  _T_872_3 = _RAND_283[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_284 = {1{`RANDOM}};
  _T_884_0 = _RAND_284[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_285 = {1{`RANDOM}};
  _T_884_1 = _RAND_285[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_286 = {1{`RANDOM}};
  _T_884_2 = _RAND_286[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_287 = {1{`RANDOM}};
  _T_884_3 = _RAND_287[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_288 = {1{`RANDOM}};
  _T_898_0 = _RAND_288[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_289 = {1{`RANDOM}};
  _T_898_1 = _RAND_289[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_290 = {1{`RANDOM}};
  _T_898_2 = _RAND_290[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_291 = {1{`RANDOM}};
  _T_898_3 = _RAND_291[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_292 = {1{`RANDOM}};
  _T_910_0 = _RAND_292[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_293 = {1{`RANDOM}};
  _T_910_1 = _RAND_293[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_294 = {1{`RANDOM}};
  _T_910_2 = _RAND_294[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_295 = {1{`RANDOM}};
  _T_910_3 = _RAND_295[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_296 = {1{`RANDOM}};
  _T_922_0 = _RAND_296[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_297 = {1{`RANDOM}};
  _T_922_1 = _RAND_297[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_298 = {1{`RANDOM}};
  _T_922_2 = _RAND_298[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_299 = {1{`RANDOM}};
  _T_922_3 = _RAND_299[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_300 = {1{`RANDOM}};
  _T_934_0 = _RAND_300[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_301 = {1{`RANDOM}};
  _T_934_1 = _RAND_301[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_302 = {1{`RANDOM}};
  _T_934_2 = _RAND_302[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_303 = {1{`RANDOM}};
  _T_934_3 = _RAND_303[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_304 = {1{`RANDOM}};
  _T_946_0 = _RAND_304[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_305 = {1{`RANDOM}};
  _T_946_1 = _RAND_305[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_306 = {1{`RANDOM}};
  _T_946_2 = _RAND_306[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_307 = {1{`RANDOM}};
  _T_946_3 = _RAND_307[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_308 = {1{`RANDOM}};
  _T_958_0 = _RAND_308[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_309 = {1{`RANDOM}};
  _T_958_1 = _RAND_309[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_310 = {1{`RANDOM}};
  _T_958_2 = _RAND_310[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_311 = {1{`RANDOM}};
  _T_958_3 = _RAND_311[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_312 = {1{`RANDOM}};
  _T_970_0 = _RAND_312[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_313 = {1{`RANDOM}};
  _T_970_1 = _RAND_313[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_314 = {1{`RANDOM}};
  _T_970_2 = _RAND_314[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_315 = {1{`RANDOM}};
  _T_970_3 = _RAND_315[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_316 = {1{`RANDOM}};
  _T_982_0 = _RAND_316[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_317 = {1{`RANDOM}};
  _T_982_1 = _RAND_317[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_318 = {1{`RANDOM}};
  _T_982_2 = _RAND_318[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_319 = {1{`RANDOM}};
  _T_982_3 = _RAND_319[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_320 = {1{`RANDOM}};
  _T_996_0 = _RAND_320[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_321 = {1{`RANDOM}};
  _T_996_1 = _RAND_321[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_322 = {1{`RANDOM}};
  _T_996_2 = _RAND_322[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_323 = {1{`RANDOM}};
  _T_996_3 = _RAND_323[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_324 = {1{`RANDOM}};
  _T_1008_0 = _RAND_324[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_325 = {1{`RANDOM}};
  _T_1008_1 = _RAND_325[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_326 = {1{`RANDOM}};
  _T_1008_2 = _RAND_326[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_327 = {1{`RANDOM}};
  _T_1008_3 = _RAND_327[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_328 = {1{`RANDOM}};
  _T_1020_0 = _RAND_328[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_329 = {1{`RANDOM}};
  _T_1020_1 = _RAND_329[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_330 = {1{`RANDOM}};
  _T_1020_2 = _RAND_330[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_331 = {1{`RANDOM}};
  _T_1020_3 = _RAND_331[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_332 = {1{`RANDOM}};
  _T_1032_0 = _RAND_332[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_333 = {1{`RANDOM}};
  _T_1032_1 = _RAND_333[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_334 = {1{`RANDOM}};
  _T_1032_2 = _RAND_334[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_335 = {1{`RANDOM}};
  _T_1032_3 = _RAND_335[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_336 = {1{`RANDOM}};
  _T_1044_0 = _RAND_336[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_337 = {1{`RANDOM}};
  _T_1044_1 = _RAND_337[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_338 = {1{`RANDOM}};
  _T_1044_2 = _RAND_338[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_339 = {1{`RANDOM}};
  _T_1044_3 = _RAND_339[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_340 = {1{`RANDOM}};
  _T_1056_0 = _RAND_340[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_341 = {1{`RANDOM}};
  _T_1056_1 = _RAND_341[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_342 = {1{`RANDOM}};
  _T_1056_2 = _RAND_342[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_343 = {1{`RANDOM}};
  _T_1056_3 = _RAND_343[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_344 = {1{`RANDOM}};
  _T_1068_0 = _RAND_344[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_345 = {1{`RANDOM}};
  _T_1068_1 = _RAND_345[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_346 = {1{`RANDOM}};
  _T_1068_2 = _RAND_346[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_347 = {1{`RANDOM}};
  _T_1068_3 = _RAND_347[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_348 = {1{`RANDOM}};
  _T_1080_0 = _RAND_348[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_349 = {1{`RANDOM}};
  _T_1080_1 = _RAND_349[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_350 = {1{`RANDOM}};
  _T_1080_2 = _RAND_350[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_351 = {1{`RANDOM}};
  _T_1080_3 = _RAND_351[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_352 = {1{`RANDOM}};
  _T_1094_0 = _RAND_352[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_353 = {1{`RANDOM}};
  _T_1094_1 = _RAND_353[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_354 = {1{`RANDOM}};
  _T_1094_2 = _RAND_354[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_355 = {1{`RANDOM}};
  _T_1094_3 = _RAND_355[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_356 = {1{`RANDOM}};
  _T_1106_0 = _RAND_356[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_357 = {1{`RANDOM}};
  _T_1106_1 = _RAND_357[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_358 = {1{`RANDOM}};
  _T_1106_2 = _RAND_358[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_359 = {1{`RANDOM}};
  _T_1106_3 = _RAND_359[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_360 = {1{`RANDOM}};
  _T_1118_0 = _RAND_360[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_361 = {1{`RANDOM}};
  _T_1118_1 = _RAND_361[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_362 = {1{`RANDOM}};
  _T_1118_2 = _RAND_362[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_363 = {1{`RANDOM}};
  _T_1118_3 = _RAND_363[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_364 = {1{`RANDOM}};
  _T_1130_0 = _RAND_364[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_365 = {1{`RANDOM}};
  _T_1130_1 = _RAND_365[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_366 = {1{`RANDOM}};
  _T_1130_2 = _RAND_366[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_367 = {1{`RANDOM}};
  _T_1130_3 = _RAND_367[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_368 = {1{`RANDOM}};
  _T_1142_0 = _RAND_368[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_369 = {1{`RANDOM}};
  _T_1142_1 = _RAND_369[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_370 = {1{`RANDOM}};
  _T_1142_2 = _RAND_370[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_371 = {1{`RANDOM}};
  _T_1142_3 = _RAND_371[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_372 = {1{`RANDOM}};
  _T_1154_0 = _RAND_372[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_373 = {1{`RANDOM}};
  _T_1154_1 = _RAND_373[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_374 = {1{`RANDOM}};
  _T_1154_2 = _RAND_374[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_375 = {1{`RANDOM}};
  _T_1154_3 = _RAND_375[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_376 = {1{`RANDOM}};
  _T_1166_0 = _RAND_376[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_377 = {1{`RANDOM}};
  _T_1166_1 = _RAND_377[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_378 = {1{`RANDOM}};
  _T_1166_2 = _RAND_378[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_379 = {1{`RANDOM}};
  _T_1166_3 = _RAND_379[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_380 = {1{`RANDOM}};
  _T_1178_0 = _RAND_380[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_381 = {1{`RANDOM}};
  _T_1178_1 = _RAND_381[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_382 = {1{`RANDOM}};
  _T_1178_2 = _RAND_382[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_383 = {1{`RANDOM}};
  _T_1178_3 = _RAND_383[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_384 = {1{`RANDOM}};
  _T_1192_0 = _RAND_384[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_385 = {1{`RANDOM}};
  _T_1192_1 = _RAND_385[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_386 = {1{`RANDOM}};
  _T_1192_2 = _RAND_386[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_387 = {1{`RANDOM}};
  _T_1192_3 = _RAND_387[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_388 = {1{`RANDOM}};
  _T_1204_0 = _RAND_388[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_389 = {1{`RANDOM}};
  _T_1204_1 = _RAND_389[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_390 = {1{`RANDOM}};
  _T_1204_2 = _RAND_390[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_391 = {1{`RANDOM}};
  _T_1204_3 = _RAND_391[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_392 = {1{`RANDOM}};
  _T_1216_0 = _RAND_392[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_393 = {1{`RANDOM}};
  _T_1216_1 = _RAND_393[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_394 = {1{`RANDOM}};
  _T_1216_2 = _RAND_394[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_395 = {1{`RANDOM}};
  _T_1216_3 = _RAND_395[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_396 = {1{`RANDOM}};
  _T_1228_0 = _RAND_396[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_397 = {1{`RANDOM}};
  _T_1228_1 = _RAND_397[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_398 = {1{`RANDOM}};
  _T_1228_2 = _RAND_398[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_399 = {1{`RANDOM}};
  _T_1228_3 = _RAND_399[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_400 = {1{`RANDOM}};
  _T_1240_0 = _RAND_400[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_401 = {1{`RANDOM}};
  _T_1240_1 = _RAND_401[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_402 = {1{`RANDOM}};
  _T_1240_2 = _RAND_402[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_403 = {1{`RANDOM}};
  _T_1240_3 = _RAND_403[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_404 = {1{`RANDOM}};
  _T_1252_0 = _RAND_404[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_405 = {1{`RANDOM}};
  _T_1252_1 = _RAND_405[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_406 = {1{`RANDOM}};
  _T_1252_2 = _RAND_406[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_407 = {1{`RANDOM}};
  _T_1252_3 = _RAND_407[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_408 = {1{`RANDOM}};
  _T_1264_0 = _RAND_408[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_409 = {1{`RANDOM}};
  _T_1264_1 = _RAND_409[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_410 = {1{`RANDOM}};
  _T_1264_2 = _RAND_410[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_411 = {1{`RANDOM}};
  _T_1264_3 = _RAND_411[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_412 = {1{`RANDOM}};
  _T_1276_0 = _RAND_412[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_413 = {1{`RANDOM}};
  _T_1276_1 = _RAND_413[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_414 = {1{`RANDOM}};
  _T_1276_2 = _RAND_414[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_415 = {1{`RANDOM}};
  _T_1276_3 = _RAND_415[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_416 = {1{`RANDOM}};
  _T_1290_0 = _RAND_416[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_417 = {1{`RANDOM}};
  _T_1290_1 = _RAND_417[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_418 = {1{`RANDOM}};
  _T_1290_2 = _RAND_418[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_419 = {1{`RANDOM}};
  _T_1290_3 = _RAND_419[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_420 = {1{`RANDOM}};
  _T_1302_0 = _RAND_420[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_421 = {1{`RANDOM}};
  _T_1302_1 = _RAND_421[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_422 = {1{`RANDOM}};
  _T_1302_2 = _RAND_422[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_423 = {1{`RANDOM}};
  _T_1302_3 = _RAND_423[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_424 = {1{`RANDOM}};
  _T_1314_0 = _RAND_424[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_425 = {1{`RANDOM}};
  _T_1314_1 = _RAND_425[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_426 = {1{`RANDOM}};
  _T_1314_2 = _RAND_426[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_427 = {1{`RANDOM}};
  _T_1314_3 = _RAND_427[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_428 = {1{`RANDOM}};
  _T_1326_0 = _RAND_428[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_429 = {1{`RANDOM}};
  _T_1326_1 = _RAND_429[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_430 = {1{`RANDOM}};
  _T_1326_2 = _RAND_430[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_431 = {1{`RANDOM}};
  _T_1326_3 = _RAND_431[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_432 = {1{`RANDOM}};
  _T_1338_0 = _RAND_432[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_433 = {1{`RANDOM}};
  _T_1338_1 = _RAND_433[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_434 = {1{`RANDOM}};
  _T_1338_2 = _RAND_434[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_435 = {1{`RANDOM}};
  _T_1338_3 = _RAND_435[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_436 = {1{`RANDOM}};
  _T_1350_0 = _RAND_436[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_437 = {1{`RANDOM}};
  _T_1350_1 = _RAND_437[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_438 = {1{`RANDOM}};
  _T_1350_2 = _RAND_438[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_439 = {1{`RANDOM}};
  _T_1350_3 = _RAND_439[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_440 = {1{`RANDOM}};
  _T_1362_0 = _RAND_440[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_441 = {1{`RANDOM}};
  _T_1362_1 = _RAND_441[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_442 = {1{`RANDOM}};
  _T_1362_2 = _RAND_442[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_443 = {1{`RANDOM}};
  _T_1362_3 = _RAND_443[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_444 = {1{`RANDOM}};
  _T_1374_0 = _RAND_444[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_445 = {1{`RANDOM}};
  _T_1374_1 = _RAND_445[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_446 = {1{`RANDOM}};
  _T_1374_2 = _RAND_446[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_447 = {1{`RANDOM}};
  _T_1374_3 = _RAND_447[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_448 = {1{`RANDOM}};
  _T_1388_0 = _RAND_448[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_449 = {1{`RANDOM}};
  _T_1388_1 = _RAND_449[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_450 = {1{`RANDOM}};
  _T_1388_2 = _RAND_450[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_451 = {1{`RANDOM}};
  _T_1388_3 = _RAND_451[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_452 = {1{`RANDOM}};
  _T_1400_0 = _RAND_452[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_453 = {1{`RANDOM}};
  _T_1400_1 = _RAND_453[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_454 = {1{`RANDOM}};
  _T_1400_2 = _RAND_454[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_455 = {1{`RANDOM}};
  _T_1400_3 = _RAND_455[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_456 = {1{`RANDOM}};
  _T_1412_0 = _RAND_456[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_457 = {1{`RANDOM}};
  _T_1412_1 = _RAND_457[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_458 = {1{`RANDOM}};
  _T_1412_2 = _RAND_458[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_459 = {1{`RANDOM}};
  _T_1412_3 = _RAND_459[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_460 = {1{`RANDOM}};
  _T_1424_0 = _RAND_460[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_461 = {1{`RANDOM}};
  _T_1424_1 = _RAND_461[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_462 = {1{`RANDOM}};
  _T_1424_2 = _RAND_462[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_463 = {1{`RANDOM}};
  _T_1424_3 = _RAND_463[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_464 = {1{`RANDOM}};
  _T_1436_0 = _RAND_464[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_465 = {1{`RANDOM}};
  _T_1436_1 = _RAND_465[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_466 = {1{`RANDOM}};
  _T_1436_2 = _RAND_466[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_467 = {1{`RANDOM}};
  _T_1436_3 = _RAND_467[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_468 = {1{`RANDOM}};
  _T_1448_0 = _RAND_468[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_469 = {1{`RANDOM}};
  _T_1448_1 = _RAND_469[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_470 = {1{`RANDOM}};
  _T_1448_2 = _RAND_470[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_471 = {1{`RANDOM}};
  _T_1448_3 = _RAND_471[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_472 = {1{`RANDOM}};
  _T_1460_0 = _RAND_472[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_473 = {1{`RANDOM}};
  _T_1460_1 = _RAND_473[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_474 = {1{`RANDOM}};
  _T_1460_2 = _RAND_474[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_475 = {1{`RANDOM}};
  _T_1460_3 = _RAND_475[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_476 = {1{`RANDOM}};
  _T_1472_0 = _RAND_476[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_477 = {1{`RANDOM}};
  _T_1472_1 = _RAND_477[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_478 = {1{`RANDOM}};
  _T_1472_2 = _RAND_478[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_479 = {1{`RANDOM}};
  _T_1472_3 = _RAND_479[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_480 = {1{`RANDOM}};
  _T_1486_0 = _RAND_480[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_481 = {1{`RANDOM}};
  _T_1486_1 = _RAND_481[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_482 = {1{`RANDOM}};
  _T_1486_2 = _RAND_482[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_483 = {1{`RANDOM}};
  _T_1486_3 = _RAND_483[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_484 = {1{`RANDOM}};
  _T_1498_0 = _RAND_484[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_485 = {1{`RANDOM}};
  _T_1498_1 = _RAND_485[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_486 = {1{`RANDOM}};
  _T_1498_2 = _RAND_486[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_487 = {1{`RANDOM}};
  _T_1498_3 = _RAND_487[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_488 = {1{`RANDOM}};
  _T_1510_0 = _RAND_488[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_489 = {1{`RANDOM}};
  _T_1510_1 = _RAND_489[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_490 = {1{`RANDOM}};
  _T_1510_2 = _RAND_490[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_491 = {1{`RANDOM}};
  _T_1510_3 = _RAND_491[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_492 = {1{`RANDOM}};
  _T_1522_0 = _RAND_492[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_493 = {1{`RANDOM}};
  _T_1522_1 = _RAND_493[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_494 = {1{`RANDOM}};
  _T_1522_2 = _RAND_494[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_495 = {1{`RANDOM}};
  _T_1522_3 = _RAND_495[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_496 = {1{`RANDOM}};
  _T_1534_0 = _RAND_496[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_497 = {1{`RANDOM}};
  _T_1534_1 = _RAND_497[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_498 = {1{`RANDOM}};
  _T_1534_2 = _RAND_498[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_499 = {1{`RANDOM}};
  _T_1534_3 = _RAND_499[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_500 = {1{`RANDOM}};
  _T_1546_0 = _RAND_500[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_501 = {1{`RANDOM}};
  _T_1546_1 = _RAND_501[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_502 = {1{`RANDOM}};
  _T_1546_2 = _RAND_502[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_503 = {1{`RANDOM}};
  _T_1546_3 = _RAND_503[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_504 = {1{`RANDOM}};
  _T_1558_0 = _RAND_504[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_505 = {1{`RANDOM}};
  _T_1558_1 = _RAND_505[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_506 = {1{`RANDOM}};
  _T_1558_2 = _RAND_506[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_507 = {1{`RANDOM}};
  _T_1558_3 = _RAND_507[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_508 = {1{`RANDOM}};
  _T_1570_0 = _RAND_508[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_509 = {1{`RANDOM}};
  _T_1570_1 = _RAND_509[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_510 = {1{`RANDOM}};
  _T_1570_2 = _RAND_510[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_511 = {1{`RANDOM}};
  _T_1570_3 = _RAND_511[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_512 = {1{`RANDOM}};
  _T_1585_0 = _RAND_512[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_513 = {1{`RANDOM}};
  _T_1585_1 = _RAND_513[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_514 = {1{`RANDOM}};
  _T_1585_2 = _RAND_514[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_515 = {1{`RANDOM}};
  _T_1594_0 = _RAND_515[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_516 = {1{`RANDOM}};
  _T_1594_1 = _RAND_516[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_517 = {1{`RANDOM}};
  _T_1594_2 = _RAND_517[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_518 = {1{`RANDOM}};
  _T_1603_0 = _RAND_518[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_519 = {1{`RANDOM}};
  _T_1603_1 = _RAND_519[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_520 = {1{`RANDOM}};
  _T_1603_2 = _RAND_520[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_521 = {1{`RANDOM}};
  _T_1612_0 = _RAND_521[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_522 = {1{`RANDOM}};
  _T_1612_1 = _RAND_522[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_523 = {1{`RANDOM}};
  _T_1612_2 = _RAND_523[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_524 = {1{`RANDOM}};
  _T_1621_0 = _RAND_524[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_525 = {1{`RANDOM}};
  _T_1621_1 = _RAND_525[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_526 = {1{`RANDOM}};
  _T_1621_2 = _RAND_526[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_527 = {1{`RANDOM}};
  _T_1630_0 = _RAND_527[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_528 = {1{`RANDOM}};
  _T_1630_1 = _RAND_528[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_529 = {1{`RANDOM}};
  _T_1630_2 = _RAND_529[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_530 = {1{`RANDOM}};
  _T_1639_0 = _RAND_530[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_531 = {1{`RANDOM}};
  _T_1639_1 = _RAND_531[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_532 = {1{`RANDOM}};
  _T_1639_2 = _RAND_532[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_533 = {1{`RANDOM}};
  _T_1648_0 = _RAND_533[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_534 = {1{`RANDOM}};
  _T_1648_1 = _RAND_534[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_535 = {1{`RANDOM}};
  _T_1648_2 = _RAND_535[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_536 = {1{`RANDOM}};
  _T_1657_0 = _RAND_536[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_537 = {1{`RANDOM}};
  _T_1657_1 = _RAND_537[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_538 = {1{`RANDOM}};
  _T_1657_2 = _RAND_538[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_539 = {1{`RANDOM}};
  _T_1666_0 = _RAND_539[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_540 = {1{`RANDOM}};
  _T_1666_1 = _RAND_540[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_541 = {1{`RANDOM}};
  _T_1666_2 = _RAND_541[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_542 = {1{`RANDOM}};
  _T_1675_0 = _RAND_542[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_543 = {1{`RANDOM}};
  _T_1675_1 = _RAND_543[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_544 = {1{`RANDOM}};
  _T_1675_2 = _RAND_544[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_545 = {1{`RANDOM}};
  _T_1684_0 = _RAND_545[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_546 = {1{`RANDOM}};
  _T_1684_1 = _RAND_546[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_547 = {1{`RANDOM}};
  _T_1684_2 = _RAND_547[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_548 = {1{`RANDOM}};
  _T_1693_0 = _RAND_548[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_549 = {1{`RANDOM}};
  _T_1693_1 = _RAND_549[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_550 = {1{`RANDOM}};
  _T_1693_2 = _RAND_550[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_551 = {1{`RANDOM}};
  _T_1702_0 = _RAND_551[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_552 = {1{`RANDOM}};
  _T_1702_1 = _RAND_552[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_553 = {1{`RANDOM}};
  _T_1702_2 = _RAND_553[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_554 = {1{`RANDOM}};
  _T_1711_0 = _RAND_554[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_555 = {1{`RANDOM}};
  _T_1711_1 = _RAND_555[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_556 = {1{`RANDOM}};
  _T_1711_2 = _RAND_556[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_557 = {1{`RANDOM}};
  _T_1720_0 = _RAND_557[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_558 = {1{`RANDOM}};
  _T_1720_1 = _RAND_558[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_559 = {1{`RANDOM}};
  _T_1720_2 = _RAND_559[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_560 = {1{`RANDOM}};
  _T_1722_0 = _RAND_560[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_561 = {1{`RANDOM}};
  _T_1722_1 = _RAND_561[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_562 = {1{`RANDOM}};
  _T_1722_2 = _RAND_562[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_563 = {1{`RANDOM}};
  _T_1722_3 = _RAND_563[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_564 = {1{`RANDOM}};
  _T_1722_4 = _RAND_564[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_565 = {1{`RANDOM}};
  _T_1722_5 = _RAND_565[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_566 = {1{`RANDOM}};
  _T_1722_6 = _RAND_566[0:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`endif // SYNTHESIS
  always @(posedge clock) begin
    if (reset) begin
      _T_16_0 <= 1'h0;
    end else begin
      _T_16_0 <= _T_9;
    end
    if (reset) begin
      _T_16_1 <= 1'h0;
    end else begin
      _T_16_1 <= _T_16_0;
    end
    if (reset) begin
      _T_16_2 <= 1'h0;
    end else begin
      _T_16_2 <= _T_16_1;
    end
    if (reset) begin
      _T_16_3 <= 1'h0;
    end else begin
      _T_16_3 <= _T_16_2;
    end
    if (reset) begin
      _T_28_0 <= 1'h0;
    end else begin
      _T_28_0 <= _T_21;
    end
    if (reset) begin
      _T_28_1 <= 1'h0;
    end else begin
      _T_28_1 <= _T_28_0;
    end
    if (reset) begin
      _T_28_2 <= 1'h0;
    end else begin
      _T_28_2 <= _T_28_1;
    end
    if (reset) begin
      _T_28_3 <= 1'h0;
    end else begin
      _T_28_3 <= _T_28_2;
    end
    if (reset) begin
      _T_40_0 <= 1'h0;
    end else begin
      _T_40_0 <= _T_33;
    end
    if (reset) begin
      _T_40_1 <= 1'h0;
    end else begin
      _T_40_1 <= _T_40_0;
    end
    if (reset) begin
      _T_40_2 <= 1'h0;
    end else begin
      _T_40_2 <= _T_40_1;
    end
    if (reset) begin
      _T_40_3 <= 1'h0;
    end else begin
      _T_40_3 <= _T_40_2;
    end
    if (reset) begin
      _T_52_0 <= 1'h0;
    end else begin
      _T_52_0 <= _T_45;
    end
    if (reset) begin
      _T_52_1 <= 1'h0;
    end else begin
      _T_52_1 <= _T_52_0;
    end
    if (reset) begin
      _T_52_2 <= 1'h0;
    end else begin
      _T_52_2 <= _T_52_1;
    end
    if (reset) begin
      _T_52_3 <= 1'h0;
    end else begin
      _T_52_3 <= _T_52_2;
    end
    if (reset) begin
      _T_64_0 <= 1'h0;
    end else begin
      _T_64_0 <= _T_57;
    end
    if (reset) begin
      _T_64_1 <= 1'h0;
    end else begin
      _T_64_1 <= _T_64_0;
    end
    if (reset) begin
      _T_64_2 <= 1'h0;
    end else begin
      _T_64_2 <= _T_64_1;
    end
    if (reset) begin
      _T_64_3 <= 1'h0;
    end else begin
      _T_64_3 <= _T_64_2;
    end
    if (reset) begin
      _T_76_0 <= 1'h0;
    end else begin
      _T_76_0 <= _T_69;
    end
    if (reset) begin
      _T_76_1 <= 1'h0;
    end else begin
      _T_76_1 <= _T_76_0;
    end
    if (reset) begin
      _T_76_2 <= 1'h0;
    end else begin
      _T_76_2 <= _T_76_1;
    end
    if (reset) begin
      _T_76_3 <= 1'h0;
    end else begin
      _T_76_3 <= _T_76_2;
    end
    if (reset) begin
      _T_88_0 <= 1'h0;
    end else begin
      _T_88_0 <= _T_81;
    end
    if (reset) begin
      _T_88_1 <= 1'h0;
    end else begin
      _T_88_1 <= _T_88_0;
    end
    if (reset) begin
      _T_88_2 <= 1'h0;
    end else begin
      _T_88_2 <= _T_88_1;
    end
    if (reset) begin
      _T_88_3 <= 1'h0;
    end else begin
      _T_88_3 <= _T_88_2;
    end
    if (reset) begin
      _T_100_0 <= 1'h0;
    end else begin
      _T_100_0 <= _T_93;
    end
    if (reset) begin
      _T_100_1 <= 1'h0;
    end else begin
      _T_100_1 <= _T_100_0;
    end
    if (reset) begin
      _T_100_2 <= 1'h0;
    end else begin
      _T_100_2 <= _T_100_1;
    end
    if (reset) begin
      _T_100_3 <= 1'h0;
    end else begin
      _T_100_3 <= _T_100_2;
    end
    if (reset) begin
      _T_114_0 <= 1'h0;
    end else begin
      _T_114_0 <= _T_21;
    end
    if (reset) begin
      _T_114_1 <= 1'h0;
    end else begin
      _T_114_1 <= _T_114_0;
    end
    if (reset) begin
      _T_114_2 <= 1'h0;
    end else begin
      _T_114_2 <= _T_114_1;
    end
    if (reset) begin
      _T_114_3 <= 1'h0;
    end else begin
      _T_114_3 <= _T_114_2;
    end
    if (reset) begin
      _T_126_0 <= 1'h0;
    end else begin
      _T_126_0 <= _T_33;
    end
    if (reset) begin
      _T_126_1 <= 1'h0;
    end else begin
      _T_126_1 <= _T_126_0;
    end
    if (reset) begin
      _T_126_2 <= 1'h0;
    end else begin
      _T_126_2 <= _T_126_1;
    end
    if (reset) begin
      _T_126_3 <= 1'h0;
    end else begin
      _T_126_3 <= _T_126_2;
    end
    if (reset) begin
      _T_138_0 <= 1'h0;
    end else begin
      _T_138_0 <= _T_45;
    end
    if (reset) begin
      _T_138_1 <= 1'h0;
    end else begin
      _T_138_1 <= _T_138_0;
    end
    if (reset) begin
      _T_138_2 <= 1'h0;
    end else begin
      _T_138_2 <= _T_138_1;
    end
    if (reset) begin
      _T_138_3 <= 1'h0;
    end else begin
      _T_138_3 <= _T_138_2;
    end
    if (reset) begin
      _T_150_0 <= 1'h0;
    end else begin
      _T_150_0 <= _T_57;
    end
    if (reset) begin
      _T_150_1 <= 1'h0;
    end else begin
      _T_150_1 <= _T_150_0;
    end
    if (reset) begin
      _T_150_2 <= 1'h0;
    end else begin
      _T_150_2 <= _T_150_1;
    end
    if (reset) begin
      _T_150_3 <= 1'h0;
    end else begin
      _T_150_3 <= _T_150_2;
    end
    if (reset) begin
      _T_162_0 <= 1'h0;
    end else begin
      _T_162_0 <= _T_69;
    end
    if (reset) begin
      _T_162_1 <= 1'h0;
    end else begin
      _T_162_1 <= _T_162_0;
    end
    if (reset) begin
      _T_162_2 <= 1'h0;
    end else begin
      _T_162_2 <= _T_162_1;
    end
    if (reset) begin
      _T_162_3 <= 1'h0;
    end else begin
      _T_162_3 <= _T_162_2;
    end
    if (reset) begin
      _T_174_0 <= 1'h0;
    end else begin
      _T_174_0 <= _T_81;
    end
    if (reset) begin
      _T_174_1 <= 1'h0;
    end else begin
      _T_174_1 <= _T_174_0;
    end
    if (reset) begin
      _T_174_2 <= 1'h0;
    end else begin
      _T_174_2 <= _T_174_1;
    end
    if (reset) begin
      _T_174_3 <= 1'h0;
    end else begin
      _T_174_3 <= _T_174_2;
    end
    if (reset) begin
      _T_186_0 <= 1'h0;
    end else begin
      _T_186_0 <= _T_93;
    end
    if (reset) begin
      _T_186_1 <= 1'h0;
    end else begin
      _T_186_1 <= _T_186_0;
    end
    if (reset) begin
      _T_186_2 <= 1'h0;
    end else begin
      _T_186_2 <= _T_186_1;
    end
    if (reset) begin
      _T_186_3 <= 1'h0;
    end else begin
      _T_186_3 <= _T_186_2;
    end
    if (reset) begin
      _T_198_0 <= 1'h0;
    end else begin
      _T_198_0 <= _T_191;
    end
    if (reset) begin
      _T_198_1 <= 1'h0;
    end else begin
      _T_198_1 <= _T_198_0;
    end
    if (reset) begin
      _T_198_2 <= 1'h0;
    end else begin
      _T_198_2 <= _T_198_1;
    end
    if (reset) begin
      _T_198_3 <= 1'h0;
    end else begin
      _T_198_3 <= _T_198_2;
    end
    if (reset) begin
      _T_212_0 <= 1'h0;
    end else begin
      _T_212_0 <= _T_33;
    end
    if (reset) begin
      _T_212_1 <= 1'h0;
    end else begin
      _T_212_1 <= _T_212_0;
    end
    if (reset) begin
      _T_212_2 <= 1'h0;
    end else begin
      _T_212_2 <= _T_212_1;
    end
    if (reset) begin
      _T_212_3 <= 1'h0;
    end else begin
      _T_212_3 <= _T_212_2;
    end
    if (reset) begin
      _T_224_0 <= 1'h0;
    end else begin
      _T_224_0 <= _T_45;
    end
    if (reset) begin
      _T_224_1 <= 1'h0;
    end else begin
      _T_224_1 <= _T_224_0;
    end
    if (reset) begin
      _T_224_2 <= 1'h0;
    end else begin
      _T_224_2 <= _T_224_1;
    end
    if (reset) begin
      _T_224_3 <= 1'h0;
    end else begin
      _T_224_3 <= _T_224_2;
    end
    if (reset) begin
      _T_236_0 <= 1'h0;
    end else begin
      _T_236_0 <= _T_57;
    end
    if (reset) begin
      _T_236_1 <= 1'h0;
    end else begin
      _T_236_1 <= _T_236_0;
    end
    if (reset) begin
      _T_236_2 <= 1'h0;
    end else begin
      _T_236_2 <= _T_236_1;
    end
    if (reset) begin
      _T_236_3 <= 1'h0;
    end else begin
      _T_236_3 <= _T_236_2;
    end
    if (reset) begin
      _T_248_0 <= 1'h0;
    end else begin
      _T_248_0 <= _T_69;
    end
    if (reset) begin
      _T_248_1 <= 1'h0;
    end else begin
      _T_248_1 <= _T_248_0;
    end
    if (reset) begin
      _T_248_2 <= 1'h0;
    end else begin
      _T_248_2 <= _T_248_1;
    end
    if (reset) begin
      _T_248_3 <= 1'h0;
    end else begin
      _T_248_3 <= _T_248_2;
    end
    if (reset) begin
      _T_260_0 <= 1'h0;
    end else begin
      _T_260_0 <= _T_81;
    end
    if (reset) begin
      _T_260_1 <= 1'h0;
    end else begin
      _T_260_1 <= _T_260_0;
    end
    if (reset) begin
      _T_260_2 <= 1'h0;
    end else begin
      _T_260_2 <= _T_260_1;
    end
    if (reset) begin
      _T_260_3 <= 1'h0;
    end else begin
      _T_260_3 <= _T_260_2;
    end
    if (reset) begin
      _T_272_0 <= 1'h0;
    end else begin
      _T_272_0 <= _T_93;
    end
    if (reset) begin
      _T_272_1 <= 1'h0;
    end else begin
      _T_272_1 <= _T_272_0;
    end
    if (reset) begin
      _T_272_2 <= 1'h0;
    end else begin
      _T_272_2 <= _T_272_1;
    end
    if (reset) begin
      _T_272_3 <= 1'h0;
    end else begin
      _T_272_3 <= _T_272_2;
    end
    if (reset) begin
      _T_284_0 <= 1'h0;
    end else begin
      _T_284_0 <= _T_191;
    end
    if (reset) begin
      _T_284_1 <= 1'h0;
    end else begin
      _T_284_1 <= _T_284_0;
    end
    if (reset) begin
      _T_284_2 <= 1'h0;
    end else begin
      _T_284_2 <= _T_284_1;
    end
    if (reset) begin
      _T_284_3 <= 1'h0;
    end else begin
      _T_284_3 <= _T_284_2;
    end
    if (reset) begin
      _T_296_0 <= 1'h0;
    end else begin
      _T_296_0 <= _T_289;
    end
    if (reset) begin
      _T_296_1 <= 1'h0;
    end else begin
      _T_296_1 <= _T_296_0;
    end
    if (reset) begin
      _T_296_2 <= 1'h0;
    end else begin
      _T_296_2 <= _T_296_1;
    end
    if (reset) begin
      _T_296_3 <= 1'h0;
    end else begin
      _T_296_3 <= _T_296_2;
    end
    if (reset) begin
      _T_310_0 <= 1'h0;
    end else begin
      _T_310_0 <= _T_45;
    end
    if (reset) begin
      _T_310_1 <= 1'h0;
    end else begin
      _T_310_1 <= _T_310_0;
    end
    if (reset) begin
      _T_310_2 <= 1'h0;
    end else begin
      _T_310_2 <= _T_310_1;
    end
    if (reset) begin
      _T_310_3 <= 1'h0;
    end else begin
      _T_310_3 <= _T_310_2;
    end
    if (reset) begin
      _T_322_0 <= 1'h0;
    end else begin
      _T_322_0 <= _T_57;
    end
    if (reset) begin
      _T_322_1 <= 1'h0;
    end else begin
      _T_322_1 <= _T_322_0;
    end
    if (reset) begin
      _T_322_2 <= 1'h0;
    end else begin
      _T_322_2 <= _T_322_1;
    end
    if (reset) begin
      _T_322_3 <= 1'h0;
    end else begin
      _T_322_3 <= _T_322_2;
    end
    if (reset) begin
      _T_334_0 <= 1'h0;
    end else begin
      _T_334_0 <= _T_69;
    end
    if (reset) begin
      _T_334_1 <= 1'h0;
    end else begin
      _T_334_1 <= _T_334_0;
    end
    if (reset) begin
      _T_334_2 <= 1'h0;
    end else begin
      _T_334_2 <= _T_334_1;
    end
    if (reset) begin
      _T_334_3 <= 1'h0;
    end else begin
      _T_334_3 <= _T_334_2;
    end
    if (reset) begin
      _T_346_0 <= 1'h0;
    end else begin
      _T_346_0 <= _T_81;
    end
    if (reset) begin
      _T_346_1 <= 1'h0;
    end else begin
      _T_346_1 <= _T_346_0;
    end
    if (reset) begin
      _T_346_2 <= 1'h0;
    end else begin
      _T_346_2 <= _T_346_1;
    end
    if (reset) begin
      _T_346_3 <= 1'h0;
    end else begin
      _T_346_3 <= _T_346_2;
    end
    if (reset) begin
      _T_358_0 <= 1'h0;
    end else begin
      _T_358_0 <= _T_93;
    end
    if (reset) begin
      _T_358_1 <= 1'h0;
    end else begin
      _T_358_1 <= _T_358_0;
    end
    if (reset) begin
      _T_358_2 <= 1'h0;
    end else begin
      _T_358_2 <= _T_358_1;
    end
    if (reset) begin
      _T_358_3 <= 1'h0;
    end else begin
      _T_358_3 <= _T_358_2;
    end
    if (reset) begin
      _T_370_0 <= 1'h0;
    end else begin
      _T_370_0 <= _T_191;
    end
    if (reset) begin
      _T_370_1 <= 1'h0;
    end else begin
      _T_370_1 <= _T_370_0;
    end
    if (reset) begin
      _T_370_2 <= 1'h0;
    end else begin
      _T_370_2 <= _T_370_1;
    end
    if (reset) begin
      _T_370_3 <= 1'h0;
    end else begin
      _T_370_3 <= _T_370_2;
    end
    if (reset) begin
      _T_382_0 <= 1'h0;
    end else begin
      _T_382_0 <= _T_289;
    end
    if (reset) begin
      _T_382_1 <= 1'h0;
    end else begin
      _T_382_1 <= _T_382_0;
    end
    if (reset) begin
      _T_382_2 <= 1'h0;
    end else begin
      _T_382_2 <= _T_382_1;
    end
    if (reset) begin
      _T_382_3 <= 1'h0;
    end else begin
      _T_382_3 <= _T_382_2;
    end
    if (reset) begin
      _T_394_0 <= 1'h0;
    end else begin
      _T_394_0 <= _T_387;
    end
    if (reset) begin
      _T_394_1 <= 1'h0;
    end else begin
      _T_394_1 <= _T_394_0;
    end
    if (reset) begin
      _T_394_2 <= 1'h0;
    end else begin
      _T_394_2 <= _T_394_1;
    end
    if (reset) begin
      _T_394_3 <= 1'h0;
    end else begin
      _T_394_3 <= _T_394_2;
    end
    if (reset) begin
      _T_408_0 <= 1'h0;
    end else begin
      _T_408_0 <= _T_57;
    end
    if (reset) begin
      _T_408_1 <= 1'h0;
    end else begin
      _T_408_1 <= _T_408_0;
    end
    if (reset) begin
      _T_408_2 <= 1'h0;
    end else begin
      _T_408_2 <= _T_408_1;
    end
    if (reset) begin
      _T_408_3 <= 1'h0;
    end else begin
      _T_408_3 <= _T_408_2;
    end
    if (reset) begin
      _T_420_0 <= 1'h0;
    end else begin
      _T_420_0 <= _T_69;
    end
    if (reset) begin
      _T_420_1 <= 1'h0;
    end else begin
      _T_420_1 <= _T_420_0;
    end
    if (reset) begin
      _T_420_2 <= 1'h0;
    end else begin
      _T_420_2 <= _T_420_1;
    end
    if (reset) begin
      _T_420_3 <= 1'h0;
    end else begin
      _T_420_3 <= _T_420_2;
    end
    if (reset) begin
      _T_432_0 <= 1'h0;
    end else begin
      _T_432_0 <= _T_81;
    end
    if (reset) begin
      _T_432_1 <= 1'h0;
    end else begin
      _T_432_1 <= _T_432_0;
    end
    if (reset) begin
      _T_432_2 <= 1'h0;
    end else begin
      _T_432_2 <= _T_432_1;
    end
    if (reset) begin
      _T_432_3 <= 1'h0;
    end else begin
      _T_432_3 <= _T_432_2;
    end
    if (reset) begin
      _T_444_0 <= 1'h0;
    end else begin
      _T_444_0 <= _T_93;
    end
    if (reset) begin
      _T_444_1 <= 1'h0;
    end else begin
      _T_444_1 <= _T_444_0;
    end
    if (reset) begin
      _T_444_2 <= 1'h0;
    end else begin
      _T_444_2 <= _T_444_1;
    end
    if (reset) begin
      _T_444_3 <= 1'h0;
    end else begin
      _T_444_3 <= _T_444_2;
    end
    if (reset) begin
      _T_456_0 <= 1'h0;
    end else begin
      _T_456_0 <= _T_191;
    end
    if (reset) begin
      _T_456_1 <= 1'h0;
    end else begin
      _T_456_1 <= _T_456_0;
    end
    if (reset) begin
      _T_456_2 <= 1'h0;
    end else begin
      _T_456_2 <= _T_456_1;
    end
    if (reset) begin
      _T_456_3 <= 1'h0;
    end else begin
      _T_456_3 <= _T_456_2;
    end
    if (reset) begin
      _T_468_0 <= 1'h0;
    end else begin
      _T_468_0 <= _T_289;
    end
    if (reset) begin
      _T_468_1 <= 1'h0;
    end else begin
      _T_468_1 <= _T_468_0;
    end
    if (reset) begin
      _T_468_2 <= 1'h0;
    end else begin
      _T_468_2 <= _T_468_1;
    end
    if (reset) begin
      _T_468_3 <= 1'h0;
    end else begin
      _T_468_3 <= _T_468_2;
    end
    if (reset) begin
      _T_480_0 <= 1'h0;
    end else begin
      _T_480_0 <= _T_387;
    end
    if (reset) begin
      _T_480_1 <= 1'h0;
    end else begin
      _T_480_1 <= _T_480_0;
    end
    if (reset) begin
      _T_480_2 <= 1'h0;
    end else begin
      _T_480_2 <= _T_480_1;
    end
    if (reset) begin
      _T_480_3 <= 1'h0;
    end else begin
      _T_480_3 <= _T_480_2;
    end
    if (reset) begin
      _T_492_0 <= 1'h0;
    end else begin
      _T_492_0 <= _T_485;
    end
    if (reset) begin
      _T_492_1 <= 1'h0;
    end else begin
      _T_492_1 <= _T_492_0;
    end
    if (reset) begin
      _T_492_2 <= 1'h0;
    end else begin
      _T_492_2 <= _T_492_1;
    end
    if (reset) begin
      _T_492_3 <= 1'h0;
    end else begin
      _T_492_3 <= _T_492_2;
    end
    if (reset) begin
      _T_506_0 <= 1'h0;
    end else begin
      _T_506_0 <= _T_69;
    end
    if (reset) begin
      _T_506_1 <= 1'h0;
    end else begin
      _T_506_1 <= _T_506_0;
    end
    if (reset) begin
      _T_506_2 <= 1'h0;
    end else begin
      _T_506_2 <= _T_506_1;
    end
    if (reset) begin
      _T_506_3 <= 1'h0;
    end else begin
      _T_506_3 <= _T_506_2;
    end
    if (reset) begin
      _T_518_0 <= 1'h0;
    end else begin
      _T_518_0 <= _T_81;
    end
    if (reset) begin
      _T_518_1 <= 1'h0;
    end else begin
      _T_518_1 <= _T_518_0;
    end
    if (reset) begin
      _T_518_2 <= 1'h0;
    end else begin
      _T_518_2 <= _T_518_1;
    end
    if (reset) begin
      _T_518_3 <= 1'h0;
    end else begin
      _T_518_3 <= _T_518_2;
    end
    if (reset) begin
      _T_530_0 <= 1'h0;
    end else begin
      _T_530_0 <= _T_93;
    end
    if (reset) begin
      _T_530_1 <= 1'h0;
    end else begin
      _T_530_1 <= _T_530_0;
    end
    if (reset) begin
      _T_530_2 <= 1'h0;
    end else begin
      _T_530_2 <= _T_530_1;
    end
    if (reset) begin
      _T_530_3 <= 1'h0;
    end else begin
      _T_530_3 <= _T_530_2;
    end
    if (reset) begin
      _T_542_0 <= 1'h0;
    end else begin
      _T_542_0 <= _T_191;
    end
    if (reset) begin
      _T_542_1 <= 1'h0;
    end else begin
      _T_542_1 <= _T_542_0;
    end
    if (reset) begin
      _T_542_2 <= 1'h0;
    end else begin
      _T_542_2 <= _T_542_1;
    end
    if (reset) begin
      _T_542_3 <= 1'h0;
    end else begin
      _T_542_3 <= _T_542_2;
    end
    if (reset) begin
      _T_554_0 <= 1'h0;
    end else begin
      _T_554_0 <= _T_289;
    end
    if (reset) begin
      _T_554_1 <= 1'h0;
    end else begin
      _T_554_1 <= _T_554_0;
    end
    if (reset) begin
      _T_554_2 <= 1'h0;
    end else begin
      _T_554_2 <= _T_554_1;
    end
    if (reset) begin
      _T_554_3 <= 1'h0;
    end else begin
      _T_554_3 <= _T_554_2;
    end
    if (reset) begin
      _T_566_0 <= 1'h0;
    end else begin
      _T_566_0 <= _T_387;
    end
    if (reset) begin
      _T_566_1 <= 1'h0;
    end else begin
      _T_566_1 <= _T_566_0;
    end
    if (reset) begin
      _T_566_2 <= 1'h0;
    end else begin
      _T_566_2 <= _T_566_1;
    end
    if (reset) begin
      _T_566_3 <= 1'h0;
    end else begin
      _T_566_3 <= _T_566_2;
    end
    if (reset) begin
      _T_578_0 <= 1'h0;
    end else begin
      _T_578_0 <= _T_485;
    end
    if (reset) begin
      _T_578_1 <= 1'h0;
    end else begin
      _T_578_1 <= _T_578_0;
    end
    if (reset) begin
      _T_578_2 <= 1'h0;
    end else begin
      _T_578_2 <= _T_578_1;
    end
    if (reset) begin
      _T_578_3 <= 1'h0;
    end else begin
      _T_578_3 <= _T_578_2;
    end
    if (reset) begin
      _T_590_0 <= 1'h0;
    end else begin
      _T_590_0 <= _T_583;
    end
    if (reset) begin
      _T_590_1 <= 1'h0;
    end else begin
      _T_590_1 <= _T_590_0;
    end
    if (reset) begin
      _T_590_2 <= 1'h0;
    end else begin
      _T_590_2 <= _T_590_1;
    end
    if (reset) begin
      _T_590_3 <= 1'h0;
    end else begin
      _T_590_3 <= _T_590_2;
    end
    if (reset) begin
      _T_604_0 <= 1'h0;
    end else begin
      _T_604_0 <= _T_81;
    end
    if (reset) begin
      _T_604_1 <= 1'h0;
    end else begin
      _T_604_1 <= _T_604_0;
    end
    if (reset) begin
      _T_604_2 <= 1'h0;
    end else begin
      _T_604_2 <= _T_604_1;
    end
    if (reset) begin
      _T_604_3 <= 1'h0;
    end else begin
      _T_604_3 <= _T_604_2;
    end
    if (reset) begin
      _T_616_0 <= 1'h0;
    end else begin
      _T_616_0 <= _T_93;
    end
    if (reset) begin
      _T_616_1 <= 1'h0;
    end else begin
      _T_616_1 <= _T_616_0;
    end
    if (reset) begin
      _T_616_2 <= 1'h0;
    end else begin
      _T_616_2 <= _T_616_1;
    end
    if (reset) begin
      _T_616_3 <= 1'h0;
    end else begin
      _T_616_3 <= _T_616_2;
    end
    if (reset) begin
      _T_628_0 <= 1'h0;
    end else begin
      _T_628_0 <= _T_191;
    end
    if (reset) begin
      _T_628_1 <= 1'h0;
    end else begin
      _T_628_1 <= _T_628_0;
    end
    if (reset) begin
      _T_628_2 <= 1'h0;
    end else begin
      _T_628_2 <= _T_628_1;
    end
    if (reset) begin
      _T_628_3 <= 1'h0;
    end else begin
      _T_628_3 <= _T_628_2;
    end
    if (reset) begin
      _T_640_0 <= 1'h0;
    end else begin
      _T_640_0 <= _T_289;
    end
    if (reset) begin
      _T_640_1 <= 1'h0;
    end else begin
      _T_640_1 <= _T_640_0;
    end
    if (reset) begin
      _T_640_2 <= 1'h0;
    end else begin
      _T_640_2 <= _T_640_1;
    end
    if (reset) begin
      _T_640_3 <= 1'h0;
    end else begin
      _T_640_3 <= _T_640_2;
    end
    if (reset) begin
      _T_652_0 <= 1'h0;
    end else begin
      _T_652_0 <= _T_387;
    end
    if (reset) begin
      _T_652_1 <= 1'h0;
    end else begin
      _T_652_1 <= _T_652_0;
    end
    if (reset) begin
      _T_652_2 <= 1'h0;
    end else begin
      _T_652_2 <= _T_652_1;
    end
    if (reset) begin
      _T_652_3 <= 1'h0;
    end else begin
      _T_652_3 <= _T_652_2;
    end
    if (reset) begin
      _T_664_0 <= 1'h0;
    end else begin
      _T_664_0 <= _T_485;
    end
    if (reset) begin
      _T_664_1 <= 1'h0;
    end else begin
      _T_664_1 <= _T_664_0;
    end
    if (reset) begin
      _T_664_2 <= 1'h0;
    end else begin
      _T_664_2 <= _T_664_1;
    end
    if (reset) begin
      _T_664_3 <= 1'h0;
    end else begin
      _T_664_3 <= _T_664_2;
    end
    if (reset) begin
      _T_676_0 <= 1'h0;
    end else begin
      _T_676_0 <= _T_583;
    end
    if (reset) begin
      _T_676_1 <= 1'h0;
    end else begin
      _T_676_1 <= _T_676_0;
    end
    if (reset) begin
      _T_676_2 <= 1'h0;
    end else begin
      _T_676_2 <= _T_676_1;
    end
    if (reset) begin
      _T_676_3 <= 1'h0;
    end else begin
      _T_676_3 <= _T_676_2;
    end
    if (reset) begin
      _T_688_0 <= 1'h0;
    end else begin
      _T_688_0 <= _T_681;
    end
    if (reset) begin
      _T_688_1 <= 1'h0;
    end else begin
      _T_688_1 <= _T_688_0;
    end
    if (reset) begin
      _T_688_2 <= 1'h0;
    end else begin
      _T_688_2 <= _T_688_1;
    end
    if (reset) begin
      _T_688_3 <= 1'h0;
    end else begin
      _T_688_3 <= _T_688_2;
    end
    if (reset) begin
      _T_702_0 <= 1'h0;
    end else begin
      _T_702_0 <= _T_93;
    end
    if (reset) begin
      _T_702_1 <= 1'h0;
    end else begin
      _T_702_1 <= _T_702_0;
    end
    if (reset) begin
      _T_702_2 <= 1'h0;
    end else begin
      _T_702_2 <= _T_702_1;
    end
    if (reset) begin
      _T_702_3 <= 1'h0;
    end else begin
      _T_702_3 <= _T_702_2;
    end
    if (reset) begin
      _T_714_0 <= 1'h0;
    end else begin
      _T_714_0 <= _T_191;
    end
    if (reset) begin
      _T_714_1 <= 1'h0;
    end else begin
      _T_714_1 <= _T_714_0;
    end
    if (reset) begin
      _T_714_2 <= 1'h0;
    end else begin
      _T_714_2 <= _T_714_1;
    end
    if (reset) begin
      _T_714_3 <= 1'h0;
    end else begin
      _T_714_3 <= _T_714_2;
    end
    if (reset) begin
      _T_726_0 <= 1'h0;
    end else begin
      _T_726_0 <= _T_289;
    end
    if (reset) begin
      _T_726_1 <= 1'h0;
    end else begin
      _T_726_1 <= _T_726_0;
    end
    if (reset) begin
      _T_726_2 <= 1'h0;
    end else begin
      _T_726_2 <= _T_726_1;
    end
    if (reset) begin
      _T_726_3 <= 1'h0;
    end else begin
      _T_726_3 <= _T_726_2;
    end
    if (reset) begin
      _T_738_0 <= 1'h0;
    end else begin
      _T_738_0 <= _T_387;
    end
    if (reset) begin
      _T_738_1 <= 1'h0;
    end else begin
      _T_738_1 <= _T_738_0;
    end
    if (reset) begin
      _T_738_2 <= 1'h0;
    end else begin
      _T_738_2 <= _T_738_1;
    end
    if (reset) begin
      _T_738_3 <= 1'h0;
    end else begin
      _T_738_3 <= _T_738_2;
    end
    if (reset) begin
      _T_750_0 <= 1'h0;
    end else begin
      _T_750_0 <= _T_485;
    end
    if (reset) begin
      _T_750_1 <= 1'h0;
    end else begin
      _T_750_1 <= _T_750_0;
    end
    if (reset) begin
      _T_750_2 <= 1'h0;
    end else begin
      _T_750_2 <= _T_750_1;
    end
    if (reset) begin
      _T_750_3 <= 1'h0;
    end else begin
      _T_750_3 <= _T_750_2;
    end
    if (reset) begin
      _T_762_0 <= 1'h0;
    end else begin
      _T_762_0 <= _T_583;
    end
    if (reset) begin
      _T_762_1 <= 1'h0;
    end else begin
      _T_762_1 <= _T_762_0;
    end
    if (reset) begin
      _T_762_2 <= 1'h0;
    end else begin
      _T_762_2 <= _T_762_1;
    end
    if (reset) begin
      _T_762_3 <= 1'h0;
    end else begin
      _T_762_3 <= _T_762_2;
    end
    if (reset) begin
      _T_774_0 <= 1'h0;
    end else begin
      _T_774_0 <= _T_681;
    end
    if (reset) begin
      _T_774_1 <= 1'h0;
    end else begin
      _T_774_1 <= _T_774_0;
    end
    if (reset) begin
      _T_774_2 <= 1'h0;
    end else begin
      _T_774_2 <= _T_774_1;
    end
    if (reset) begin
      _T_774_3 <= 1'h0;
    end else begin
      _T_774_3 <= _T_774_2;
    end
    if (reset) begin
      _T_786_0 <= 1'h0;
    end else begin
      _T_786_0 <= _T_779;
    end
    if (reset) begin
      _T_786_1 <= 1'h0;
    end else begin
      _T_786_1 <= _T_786_0;
    end
    if (reset) begin
      _T_786_2 <= 1'h0;
    end else begin
      _T_786_2 <= _T_786_1;
    end
    if (reset) begin
      _T_786_3 <= 1'h0;
    end else begin
      _T_786_3 <= _T_786_2;
    end
    if (reset) begin
      _T_800_0 <= 1'h0;
    end else begin
      _T_800_0 <= _T_191;
    end
    if (reset) begin
      _T_800_1 <= 1'h0;
    end else begin
      _T_800_1 <= _T_800_0;
    end
    if (reset) begin
      _T_800_2 <= 1'h0;
    end else begin
      _T_800_2 <= _T_800_1;
    end
    if (reset) begin
      _T_800_3 <= 1'h0;
    end else begin
      _T_800_3 <= _T_800_2;
    end
    if (reset) begin
      _T_812_0 <= 1'h0;
    end else begin
      _T_812_0 <= _T_289;
    end
    if (reset) begin
      _T_812_1 <= 1'h0;
    end else begin
      _T_812_1 <= _T_812_0;
    end
    if (reset) begin
      _T_812_2 <= 1'h0;
    end else begin
      _T_812_2 <= _T_812_1;
    end
    if (reset) begin
      _T_812_3 <= 1'h0;
    end else begin
      _T_812_3 <= _T_812_2;
    end
    if (reset) begin
      _T_824_0 <= 1'h0;
    end else begin
      _T_824_0 <= _T_387;
    end
    if (reset) begin
      _T_824_1 <= 1'h0;
    end else begin
      _T_824_1 <= _T_824_0;
    end
    if (reset) begin
      _T_824_2 <= 1'h0;
    end else begin
      _T_824_2 <= _T_824_1;
    end
    if (reset) begin
      _T_824_3 <= 1'h0;
    end else begin
      _T_824_3 <= _T_824_2;
    end
    if (reset) begin
      _T_836_0 <= 1'h0;
    end else begin
      _T_836_0 <= _T_485;
    end
    if (reset) begin
      _T_836_1 <= 1'h0;
    end else begin
      _T_836_1 <= _T_836_0;
    end
    if (reset) begin
      _T_836_2 <= 1'h0;
    end else begin
      _T_836_2 <= _T_836_1;
    end
    if (reset) begin
      _T_836_3 <= 1'h0;
    end else begin
      _T_836_3 <= _T_836_2;
    end
    if (reset) begin
      _T_848_0 <= 1'h0;
    end else begin
      _T_848_0 <= _T_583;
    end
    if (reset) begin
      _T_848_1 <= 1'h0;
    end else begin
      _T_848_1 <= _T_848_0;
    end
    if (reset) begin
      _T_848_2 <= 1'h0;
    end else begin
      _T_848_2 <= _T_848_1;
    end
    if (reset) begin
      _T_848_3 <= 1'h0;
    end else begin
      _T_848_3 <= _T_848_2;
    end
    if (reset) begin
      _T_860_0 <= 1'h0;
    end else begin
      _T_860_0 <= _T_681;
    end
    if (reset) begin
      _T_860_1 <= 1'h0;
    end else begin
      _T_860_1 <= _T_860_0;
    end
    if (reset) begin
      _T_860_2 <= 1'h0;
    end else begin
      _T_860_2 <= _T_860_1;
    end
    if (reset) begin
      _T_860_3 <= 1'h0;
    end else begin
      _T_860_3 <= _T_860_2;
    end
    if (reset) begin
      _T_872_0 <= 1'h0;
    end else begin
      _T_872_0 <= _T_779;
    end
    if (reset) begin
      _T_872_1 <= 1'h0;
    end else begin
      _T_872_1 <= _T_872_0;
    end
    if (reset) begin
      _T_872_2 <= 1'h0;
    end else begin
      _T_872_2 <= _T_872_1;
    end
    if (reset) begin
      _T_872_3 <= 1'h0;
    end else begin
      _T_872_3 <= _T_872_2;
    end
    if (reset) begin
      _T_884_0 <= 1'h0;
    end else begin
      _T_884_0 <= _T_877;
    end
    if (reset) begin
      _T_884_1 <= 1'h0;
    end else begin
      _T_884_1 <= _T_884_0;
    end
    if (reset) begin
      _T_884_2 <= 1'h0;
    end else begin
      _T_884_2 <= _T_884_1;
    end
    if (reset) begin
      _T_884_3 <= 1'h0;
    end else begin
      _T_884_3 <= _T_884_2;
    end
    if (reset) begin
      _T_898_0 <= 1'h0;
    end else begin
      _T_898_0 <= _T_289;
    end
    if (reset) begin
      _T_898_1 <= 1'h0;
    end else begin
      _T_898_1 <= _T_898_0;
    end
    if (reset) begin
      _T_898_2 <= 1'h0;
    end else begin
      _T_898_2 <= _T_898_1;
    end
    if (reset) begin
      _T_898_3 <= 1'h0;
    end else begin
      _T_898_3 <= _T_898_2;
    end
    if (reset) begin
      _T_910_0 <= 1'h0;
    end else begin
      _T_910_0 <= _T_387;
    end
    if (reset) begin
      _T_910_1 <= 1'h0;
    end else begin
      _T_910_1 <= _T_910_0;
    end
    if (reset) begin
      _T_910_2 <= 1'h0;
    end else begin
      _T_910_2 <= _T_910_1;
    end
    if (reset) begin
      _T_910_3 <= 1'h0;
    end else begin
      _T_910_3 <= _T_910_2;
    end
    if (reset) begin
      _T_922_0 <= 1'h0;
    end else begin
      _T_922_0 <= _T_485;
    end
    if (reset) begin
      _T_922_1 <= 1'h0;
    end else begin
      _T_922_1 <= _T_922_0;
    end
    if (reset) begin
      _T_922_2 <= 1'h0;
    end else begin
      _T_922_2 <= _T_922_1;
    end
    if (reset) begin
      _T_922_3 <= 1'h0;
    end else begin
      _T_922_3 <= _T_922_2;
    end
    if (reset) begin
      _T_934_0 <= 1'h0;
    end else begin
      _T_934_0 <= _T_583;
    end
    if (reset) begin
      _T_934_1 <= 1'h0;
    end else begin
      _T_934_1 <= _T_934_0;
    end
    if (reset) begin
      _T_934_2 <= 1'h0;
    end else begin
      _T_934_2 <= _T_934_1;
    end
    if (reset) begin
      _T_934_3 <= 1'h0;
    end else begin
      _T_934_3 <= _T_934_2;
    end
    if (reset) begin
      _T_946_0 <= 1'h0;
    end else begin
      _T_946_0 <= _T_681;
    end
    if (reset) begin
      _T_946_1 <= 1'h0;
    end else begin
      _T_946_1 <= _T_946_0;
    end
    if (reset) begin
      _T_946_2 <= 1'h0;
    end else begin
      _T_946_2 <= _T_946_1;
    end
    if (reset) begin
      _T_946_3 <= 1'h0;
    end else begin
      _T_946_3 <= _T_946_2;
    end
    if (reset) begin
      _T_958_0 <= 1'h0;
    end else begin
      _T_958_0 <= _T_779;
    end
    if (reset) begin
      _T_958_1 <= 1'h0;
    end else begin
      _T_958_1 <= _T_958_0;
    end
    if (reset) begin
      _T_958_2 <= 1'h0;
    end else begin
      _T_958_2 <= _T_958_1;
    end
    if (reset) begin
      _T_958_3 <= 1'h0;
    end else begin
      _T_958_3 <= _T_958_2;
    end
    if (reset) begin
      _T_970_0 <= 1'h0;
    end else begin
      _T_970_0 <= _T_877;
    end
    if (reset) begin
      _T_970_1 <= 1'h0;
    end else begin
      _T_970_1 <= _T_970_0;
    end
    if (reset) begin
      _T_970_2 <= 1'h0;
    end else begin
      _T_970_2 <= _T_970_1;
    end
    if (reset) begin
      _T_970_3 <= 1'h0;
    end else begin
      _T_970_3 <= _T_970_2;
    end
    if (reset) begin
      _T_982_0 <= 1'h0;
    end else begin
      _T_982_0 <= _T_975;
    end
    if (reset) begin
      _T_982_1 <= 1'h0;
    end else begin
      _T_982_1 <= _T_982_0;
    end
    if (reset) begin
      _T_982_2 <= 1'h0;
    end else begin
      _T_982_2 <= _T_982_1;
    end
    if (reset) begin
      _T_982_3 <= 1'h0;
    end else begin
      _T_982_3 <= _T_982_2;
    end
    if (reset) begin
      _T_996_0 <= 1'h0;
    end else begin
      _T_996_0 <= _T_387;
    end
    if (reset) begin
      _T_996_1 <= 1'h0;
    end else begin
      _T_996_1 <= _T_996_0;
    end
    if (reset) begin
      _T_996_2 <= 1'h0;
    end else begin
      _T_996_2 <= _T_996_1;
    end
    if (reset) begin
      _T_996_3 <= 1'h0;
    end else begin
      _T_996_3 <= _T_996_2;
    end
    if (reset) begin
      _T_1008_0 <= 1'h0;
    end else begin
      _T_1008_0 <= _T_485;
    end
    if (reset) begin
      _T_1008_1 <= 1'h0;
    end else begin
      _T_1008_1 <= _T_1008_0;
    end
    if (reset) begin
      _T_1008_2 <= 1'h0;
    end else begin
      _T_1008_2 <= _T_1008_1;
    end
    if (reset) begin
      _T_1008_3 <= 1'h0;
    end else begin
      _T_1008_3 <= _T_1008_2;
    end
    if (reset) begin
      _T_1020_0 <= 1'h0;
    end else begin
      _T_1020_0 <= _T_583;
    end
    if (reset) begin
      _T_1020_1 <= 1'h0;
    end else begin
      _T_1020_1 <= _T_1020_0;
    end
    if (reset) begin
      _T_1020_2 <= 1'h0;
    end else begin
      _T_1020_2 <= _T_1020_1;
    end
    if (reset) begin
      _T_1020_3 <= 1'h0;
    end else begin
      _T_1020_3 <= _T_1020_2;
    end
    if (reset) begin
      _T_1032_0 <= 1'h0;
    end else begin
      _T_1032_0 <= _T_681;
    end
    if (reset) begin
      _T_1032_1 <= 1'h0;
    end else begin
      _T_1032_1 <= _T_1032_0;
    end
    if (reset) begin
      _T_1032_2 <= 1'h0;
    end else begin
      _T_1032_2 <= _T_1032_1;
    end
    if (reset) begin
      _T_1032_3 <= 1'h0;
    end else begin
      _T_1032_3 <= _T_1032_2;
    end
    if (reset) begin
      _T_1044_0 <= 1'h0;
    end else begin
      _T_1044_0 <= _T_779;
    end
    if (reset) begin
      _T_1044_1 <= 1'h0;
    end else begin
      _T_1044_1 <= _T_1044_0;
    end
    if (reset) begin
      _T_1044_2 <= 1'h0;
    end else begin
      _T_1044_2 <= _T_1044_1;
    end
    if (reset) begin
      _T_1044_3 <= 1'h0;
    end else begin
      _T_1044_3 <= _T_1044_2;
    end
    if (reset) begin
      _T_1056_0 <= 1'h0;
    end else begin
      _T_1056_0 <= _T_877;
    end
    if (reset) begin
      _T_1056_1 <= 1'h0;
    end else begin
      _T_1056_1 <= _T_1056_0;
    end
    if (reset) begin
      _T_1056_2 <= 1'h0;
    end else begin
      _T_1056_2 <= _T_1056_1;
    end
    if (reset) begin
      _T_1056_3 <= 1'h0;
    end else begin
      _T_1056_3 <= _T_1056_2;
    end
    if (reset) begin
      _T_1068_0 <= 1'h0;
    end else begin
      _T_1068_0 <= _T_975;
    end
    if (reset) begin
      _T_1068_1 <= 1'h0;
    end else begin
      _T_1068_1 <= _T_1068_0;
    end
    if (reset) begin
      _T_1068_2 <= 1'h0;
    end else begin
      _T_1068_2 <= _T_1068_1;
    end
    if (reset) begin
      _T_1068_3 <= 1'h0;
    end else begin
      _T_1068_3 <= _T_1068_2;
    end
    if (reset) begin
      _T_1080_0 <= 1'h0;
    end else begin
      _T_1080_0 <= _T_1073;
    end
    if (reset) begin
      _T_1080_1 <= 1'h0;
    end else begin
      _T_1080_1 <= _T_1080_0;
    end
    if (reset) begin
      _T_1080_2 <= 1'h0;
    end else begin
      _T_1080_2 <= _T_1080_1;
    end
    if (reset) begin
      _T_1080_3 <= 1'h0;
    end else begin
      _T_1080_3 <= _T_1080_2;
    end
    if (reset) begin
      _T_1094_0 <= 1'h0;
    end else begin
      _T_1094_0 <= _T_485;
    end
    if (reset) begin
      _T_1094_1 <= 1'h0;
    end else begin
      _T_1094_1 <= _T_1094_0;
    end
    if (reset) begin
      _T_1094_2 <= 1'h0;
    end else begin
      _T_1094_2 <= _T_1094_1;
    end
    if (reset) begin
      _T_1094_3 <= 1'h0;
    end else begin
      _T_1094_3 <= _T_1094_2;
    end
    if (reset) begin
      _T_1106_0 <= 1'h0;
    end else begin
      _T_1106_0 <= _T_583;
    end
    if (reset) begin
      _T_1106_1 <= 1'h0;
    end else begin
      _T_1106_1 <= _T_1106_0;
    end
    if (reset) begin
      _T_1106_2 <= 1'h0;
    end else begin
      _T_1106_2 <= _T_1106_1;
    end
    if (reset) begin
      _T_1106_3 <= 1'h0;
    end else begin
      _T_1106_3 <= _T_1106_2;
    end
    if (reset) begin
      _T_1118_0 <= 1'h0;
    end else begin
      _T_1118_0 <= _T_681;
    end
    if (reset) begin
      _T_1118_1 <= 1'h0;
    end else begin
      _T_1118_1 <= _T_1118_0;
    end
    if (reset) begin
      _T_1118_2 <= 1'h0;
    end else begin
      _T_1118_2 <= _T_1118_1;
    end
    if (reset) begin
      _T_1118_3 <= 1'h0;
    end else begin
      _T_1118_3 <= _T_1118_2;
    end
    if (reset) begin
      _T_1130_0 <= 1'h0;
    end else begin
      _T_1130_0 <= _T_779;
    end
    if (reset) begin
      _T_1130_1 <= 1'h0;
    end else begin
      _T_1130_1 <= _T_1130_0;
    end
    if (reset) begin
      _T_1130_2 <= 1'h0;
    end else begin
      _T_1130_2 <= _T_1130_1;
    end
    if (reset) begin
      _T_1130_3 <= 1'h0;
    end else begin
      _T_1130_3 <= _T_1130_2;
    end
    if (reset) begin
      _T_1142_0 <= 1'h0;
    end else begin
      _T_1142_0 <= _T_877;
    end
    if (reset) begin
      _T_1142_1 <= 1'h0;
    end else begin
      _T_1142_1 <= _T_1142_0;
    end
    if (reset) begin
      _T_1142_2 <= 1'h0;
    end else begin
      _T_1142_2 <= _T_1142_1;
    end
    if (reset) begin
      _T_1142_3 <= 1'h0;
    end else begin
      _T_1142_3 <= _T_1142_2;
    end
    if (reset) begin
      _T_1154_0 <= 1'h0;
    end else begin
      _T_1154_0 <= _T_975;
    end
    if (reset) begin
      _T_1154_1 <= 1'h0;
    end else begin
      _T_1154_1 <= _T_1154_0;
    end
    if (reset) begin
      _T_1154_2 <= 1'h0;
    end else begin
      _T_1154_2 <= _T_1154_1;
    end
    if (reset) begin
      _T_1154_3 <= 1'h0;
    end else begin
      _T_1154_3 <= _T_1154_2;
    end
    if (reset) begin
      _T_1166_0 <= 1'h0;
    end else begin
      _T_1166_0 <= _T_1073;
    end
    if (reset) begin
      _T_1166_1 <= 1'h0;
    end else begin
      _T_1166_1 <= _T_1166_0;
    end
    if (reset) begin
      _T_1166_2 <= 1'h0;
    end else begin
      _T_1166_2 <= _T_1166_1;
    end
    if (reset) begin
      _T_1166_3 <= 1'h0;
    end else begin
      _T_1166_3 <= _T_1166_2;
    end
    if (reset) begin
      _T_1178_0 <= 1'h0;
    end else begin
      _T_1178_0 <= _T_1171;
    end
    if (reset) begin
      _T_1178_1 <= 1'h0;
    end else begin
      _T_1178_1 <= _T_1178_0;
    end
    if (reset) begin
      _T_1178_2 <= 1'h0;
    end else begin
      _T_1178_2 <= _T_1178_1;
    end
    if (reset) begin
      _T_1178_3 <= 1'h0;
    end else begin
      _T_1178_3 <= _T_1178_2;
    end
    if (reset) begin
      _T_1192_0 <= 1'h0;
    end else begin
      _T_1192_0 <= _T_583;
    end
    if (reset) begin
      _T_1192_1 <= 1'h0;
    end else begin
      _T_1192_1 <= _T_1192_0;
    end
    if (reset) begin
      _T_1192_2 <= 1'h0;
    end else begin
      _T_1192_2 <= _T_1192_1;
    end
    if (reset) begin
      _T_1192_3 <= 1'h0;
    end else begin
      _T_1192_3 <= _T_1192_2;
    end
    if (reset) begin
      _T_1204_0 <= 1'h0;
    end else begin
      _T_1204_0 <= _T_681;
    end
    if (reset) begin
      _T_1204_1 <= 1'h0;
    end else begin
      _T_1204_1 <= _T_1204_0;
    end
    if (reset) begin
      _T_1204_2 <= 1'h0;
    end else begin
      _T_1204_2 <= _T_1204_1;
    end
    if (reset) begin
      _T_1204_3 <= 1'h0;
    end else begin
      _T_1204_3 <= _T_1204_2;
    end
    if (reset) begin
      _T_1216_0 <= 1'h0;
    end else begin
      _T_1216_0 <= _T_779;
    end
    if (reset) begin
      _T_1216_1 <= 1'h0;
    end else begin
      _T_1216_1 <= _T_1216_0;
    end
    if (reset) begin
      _T_1216_2 <= 1'h0;
    end else begin
      _T_1216_2 <= _T_1216_1;
    end
    if (reset) begin
      _T_1216_3 <= 1'h0;
    end else begin
      _T_1216_3 <= _T_1216_2;
    end
    if (reset) begin
      _T_1228_0 <= 1'h0;
    end else begin
      _T_1228_0 <= _T_877;
    end
    if (reset) begin
      _T_1228_1 <= 1'h0;
    end else begin
      _T_1228_1 <= _T_1228_0;
    end
    if (reset) begin
      _T_1228_2 <= 1'h0;
    end else begin
      _T_1228_2 <= _T_1228_1;
    end
    if (reset) begin
      _T_1228_3 <= 1'h0;
    end else begin
      _T_1228_3 <= _T_1228_2;
    end
    if (reset) begin
      _T_1240_0 <= 1'h0;
    end else begin
      _T_1240_0 <= _T_975;
    end
    if (reset) begin
      _T_1240_1 <= 1'h0;
    end else begin
      _T_1240_1 <= _T_1240_0;
    end
    if (reset) begin
      _T_1240_2 <= 1'h0;
    end else begin
      _T_1240_2 <= _T_1240_1;
    end
    if (reset) begin
      _T_1240_3 <= 1'h0;
    end else begin
      _T_1240_3 <= _T_1240_2;
    end
    if (reset) begin
      _T_1252_0 <= 1'h0;
    end else begin
      _T_1252_0 <= _T_1073;
    end
    if (reset) begin
      _T_1252_1 <= 1'h0;
    end else begin
      _T_1252_1 <= _T_1252_0;
    end
    if (reset) begin
      _T_1252_2 <= 1'h0;
    end else begin
      _T_1252_2 <= _T_1252_1;
    end
    if (reset) begin
      _T_1252_3 <= 1'h0;
    end else begin
      _T_1252_3 <= _T_1252_2;
    end
    if (reset) begin
      _T_1264_0 <= 1'h0;
    end else begin
      _T_1264_0 <= _T_1171;
    end
    if (reset) begin
      _T_1264_1 <= 1'h0;
    end else begin
      _T_1264_1 <= _T_1264_0;
    end
    if (reset) begin
      _T_1264_2 <= 1'h0;
    end else begin
      _T_1264_2 <= _T_1264_1;
    end
    if (reset) begin
      _T_1264_3 <= 1'h0;
    end else begin
      _T_1264_3 <= _T_1264_2;
    end
    if (reset) begin
      _T_1276_0 <= 1'h0;
    end else begin
      _T_1276_0 <= _T_1269;
    end
    if (reset) begin
      _T_1276_1 <= 1'h0;
    end else begin
      _T_1276_1 <= _T_1276_0;
    end
    if (reset) begin
      _T_1276_2 <= 1'h0;
    end else begin
      _T_1276_2 <= _T_1276_1;
    end
    if (reset) begin
      _T_1276_3 <= 1'h0;
    end else begin
      _T_1276_3 <= _T_1276_2;
    end
    if (reset) begin
      _T_1290_0 <= 1'h0;
    end else begin
      _T_1290_0 <= _T_681;
    end
    if (reset) begin
      _T_1290_1 <= 1'h0;
    end else begin
      _T_1290_1 <= _T_1290_0;
    end
    if (reset) begin
      _T_1290_2 <= 1'h0;
    end else begin
      _T_1290_2 <= _T_1290_1;
    end
    if (reset) begin
      _T_1290_3 <= 1'h0;
    end else begin
      _T_1290_3 <= _T_1290_2;
    end
    if (reset) begin
      _T_1302_0 <= 1'h0;
    end else begin
      _T_1302_0 <= _T_779;
    end
    if (reset) begin
      _T_1302_1 <= 1'h0;
    end else begin
      _T_1302_1 <= _T_1302_0;
    end
    if (reset) begin
      _T_1302_2 <= 1'h0;
    end else begin
      _T_1302_2 <= _T_1302_1;
    end
    if (reset) begin
      _T_1302_3 <= 1'h0;
    end else begin
      _T_1302_3 <= _T_1302_2;
    end
    if (reset) begin
      _T_1314_0 <= 1'h0;
    end else begin
      _T_1314_0 <= _T_877;
    end
    if (reset) begin
      _T_1314_1 <= 1'h0;
    end else begin
      _T_1314_1 <= _T_1314_0;
    end
    if (reset) begin
      _T_1314_2 <= 1'h0;
    end else begin
      _T_1314_2 <= _T_1314_1;
    end
    if (reset) begin
      _T_1314_3 <= 1'h0;
    end else begin
      _T_1314_3 <= _T_1314_2;
    end
    if (reset) begin
      _T_1326_0 <= 1'h0;
    end else begin
      _T_1326_0 <= _T_975;
    end
    if (reset) begin
      _T_1326_1 <= 1'h0;
    end else begin
      _T_1326_1 <= _T_1326_0;
    end
    if (reset) begin
      _T_1326_2 <= 1'h0;
    end else begin
      _T_1326_2 <= _T_1326_1;
    end
    if (reset) begin
      _T_1326_3 <= 1'h0;
    end else begin
      _T_1326_3 <= _T_1326_2;
    end
    if (reset) begin
      _T_1338_0 <= 1'h0;
    end else begin
      _T_1338_0 <= _T_1073;
    end
    if (reset) begin
      _T_1338_1 <= 1'h0;
    end else begin
      _T_1338_1 <= _T_1338_0;
    end
    if (reset) begin
      _T_1338_2 <= 1'h0;
    end else begin
      _T_1338_2 <= _T_1338_1;
    end
    if (reset) begin
      _T_1338_3 <= 1'h0;
    end else begin
      _T_1338_3 <= _T_1338_2;
    end
    if (reset) begin
      _T_1350_0 <= 1'h0;
    end else begin
      _T_1350_0 <= _T_1171;
    end
    if (reset) begin
      _T_1350_1 <= 1'h0;
    end else begin
      _T_1350_1 <= _T_1350_0;
    end
    if (reset) begin
      _T_1350_2 <= 1'h0;
    end else begin
      _T_1350_2 <= _T_1350_1;
    end
    if (reset) begin
      _T_1350_3 <= 1'h0;
    end else begin
      _T_1350_3 <= _T_1350_2;
    end
    if (reset) begin
      _T_1362_0 <= 1'h0;
    end else begin
      _T_1362_0 <= _T_1269;
    end
    if (reset) begin
      _T_1362_1 <= 1'h0;
    end else begin
      _T_1362_1 <= _T_1362_0;
    end
    if (reset) begin
      _T_1362_2 <= 1'h0;
    end else begin
      _T_1362_2 <= _T_1362_1;
    end
    if (reset) begin
      _T_1362_3 <= 1'h0;
    end else begin
      _T_1362_3 <= _T_1362_2;
    end
    if (reset) begin
      _T_1374_0 <= 1'h0;
    end else begin
      _T_1374_0 <= _T_1367;
    end
    if (reset) begin
      _T_1374_1 <= 1'h0;
    end else begin
      _T_1374_1 <= _T_1374_0;
    end
    if (reset) begin
      _T_1374_2 <= 1'h0;
    end else begin
      _T_1374_2 <= _T_1374_1;
    end
    if (reset) begin
      _T_1374_3 <= 1'h0;
    end else begin
      _T_1374_3 <= _T_1374_2;
    end
    if (reset) begin
      _T_1388_0 <= 1'h0;
    end else begin
      _T_1388_0 <= _T_779;
    end
    if (reset) begin
      _T_1388_1 <= 1'h0;
    end else begin
      _T_1388_1 <= _T_1388_0;
    end
    if (reset) begin
      _T_1388_2 <= 1'h0;
    end else begin
      _T_1388_2 <= _T_1388_1;
    end
    if (reset) begin
      _T_1388_3 <= 1'h0;
    end else begin
      _T_1388_3 <= _T_1388_2;
    end
    if (reset) begin
      _T_1400_0 <= 1'h0;
    end else begin
      _T_1400_0 <= _T_877;
    end
    if (reset) begin
      _T_1400_1 <= 1'h0;
    end else begin
      _T_1400_1 <= _T_1400_0;
    end
    if (reset) begin
      _T_1400_2 <= 1'h0;
    end else begin
      _T_1400_2 <= _T_1400_1;
    end
    if (reset) begin
      _T_1400_3 <= 1'h0;
    end else begin
      _T_1400_3 <= _T_1400_2;
    end
    if (reset) begin
      _T_1412_0 <= 1'h0;
    end else begin
      _T_1412_0 <= _T_975;
    end
    if (reset) begin
      _T_1412_1 <= 1'h0;
    end else begin
      _T_1412_1 <= _T_1412_0;
    end
    if (reset) begin
      _T_1412_2 <= 1'h0;
    end else begin
      _T_1412_2 <= _T_1412_1;
    end
    if (reset) begin
      _T_1412_3 <= 1'h0;
    end else begin
      _T_1412_3 <= _T_1412_2;
    end
    if (reset) begin
      _T_1424_0 <= 1'h0;
    end else begin
      _T_1424_0 <= _T_1073;
    end
    if (reset) begin
      _T_1424_1 <= 1'h0;
    end else begin
      _T_1424_1 <= _T_1424_0;
    end
    if (reset) begin
      _T_1424_2 <= 1'h0;
    end else begin
      _T_1424_2 <= _T_1424_1;
    end
    if (reset) begin
      _T_1424_3 <= 1'h0;
    end else begin
      _T_1424_3 <= _T_1424_2;
    end
    if (reset) begin
      _T_1436_0 <= 1'h0;
    end else begin
      _T_1436_0 <= _T_1171;
    end
    if (reset) begin
      _T_1436_1 <= 1'h0;
    end else begin
      _T_1436_1 <= _T_1436_0;
    end
    if (reset) begin
      _T_1436_2 <= 1'h0;
    end else begin
      _T_1436_2 <= _T_1436_1;
    end
    if (reset) begin
      _T_1436_3 <= 1'h0;
    end else begin
      _T_1436_3 <= _T_1436_2;
    end
    if (reset) begin
      _T_1448_0 <= 1'h0;
    end else begin
      _T_1448_0 <= _T_1269;
    end
    if (reset) begin
      _T_1448_1 <= 1'h0;
    end else begin
      _T_1448_1 <= _T_1448_0;
    end
    if (reset) begin
      _T_1448_2 <= 1'h0;
    end else begin
      _T_1448_2 <= _T_1448_1;
    end
    if (reset) begin
      _T_1448_3 <= 1'h0;
    end else begin
      _T_1448_3 <= _T_1448_2;
    end
    if (reset) begin
      _T_1460_0 <= 1'h0;
    end else begin
      _T_1460_0 <= _T_1367;
    end
    if (reset) begin
      _T_1460_1 <= 1'h0;
    end else begin
      _T_1460_1 <= _T_1460_0;
    end
    if (reset) begin
      _T_1460_2 <= 1'h0;
    end else begin
      _T_1460_2 <= _T_1460_1;
    end
    if (reset) begin
      _T_1460_3 <= 1'h0;
    end else begin
      _T_1460_3 <= _T_1460_2;
    end
    if (reset) begin
      _T_1472_0 <= 1'h0;
    end else begin
      _T_1472_0 <= _T_1465;
    end
    if (reset) begin
      _T_1472_1 <= 1'h0;
    end else begin
      _T_1472_1 <= _T_1472_0;
    end
    if (reset) begin
      _T_1472_2 <= 1'h0;
    end else begin
      _T_1472_2 <= _T_1472_1;
    end
    if (reset) begin
      _T_1472_3 <= 1'h0;
    end else begin
      _T_1472_3 <= _T_1472_2;
    end
    if (reset) begin
      _T_1486_0 <= 1'h0;
    end else begin
      _T_1486_0 <= _T_877;
    end
    if (reset) begin
      _T_1486_1 <= 1'h0;
    end else begin
      _T_1486_1 <= _T_1486_0;
    end
    if (reset) begin
      _T_1486_2 <= 1'h0;
    end else begin
      _T_1486_2 <= _T_1486_1;
    end
    if (reset) begin
      _T_1486_3 <= 1'h0;
    end else begin
      _T_1486_3 <= _T_1486_2;
    end
    if (reset) begin
      _T_1498_0 <= 1'h0;
    end else begin
      _T_1498_0 <= _T_975;
    end
    if (reset) begin
      _T_1498_1 <= 1'h0;
    end else begin
      _T_1498_1 <= _T_1498_0;
    end
    if (reset) begin
      _T_1498_2 <= 1'h0;
    end else begin
      _T_1498_2 <= _T_1498_1;
    end
    if (reset) begin
      _T_1498_3 <= 1'h0;
    end else begin
      _T_1498_3 <= _T_1498_2;
    end
    if (reset) begin
      _T_1510_0 <= 1'h0;
    end else begin
      _T_1510_0 <= _T_1073;
    end
    if (reset) begin
      _T_1510_1 <= 1'h0;
    end else begin
      _T_1510_1 <= _T_1510_0;
    end
    if (reset) begin
      _T_1510_2 <= 1'h0;
    end else begin
      _T_1510_2 <= _T_1510_1;
    end
    if (reset) begin
      _T_1510_3 <= 1'h0;
    end else begin
      _T_1510_3 <= _T_1510_2;
    end
    if (reset) begin
      _T_1522_0 <= 1'h0;
    end else begin
      _T_1522_0 <= _T_1171;
    end
    if (reset) begin
      _T_1522_1 <= 1'h0;
    end else begin
      _T_1522_1 <= _T_1522_0;
    end
    if (reset) begin
      _T_1522_2 <= 1'h0;
    end else begin
      _T_1522_2 <= _T_1522_1;
    end
    if (reset) begin
      _T_1522_3 <= 1'h0;
    end else begin
      _T_1522_3 <= _T_1522_2;
    end
    if (reset) begin
      _T_1534_0 <= 1'h0;
    end else begin
      _T_1534_0 <= _T_1269;
    end
    if (reset) begin
      _T_1534_1 <= 1'h0;
    end else begin
      _T_1534_1 <= _T_1534_0;
    end
    if (reset) begin
      _T_1534_2 <= 1'h0;
    end else begin
      _T_1534_2 <= _T_1534_1;
    end
    if (reset) begin
      _T_1534_3 <= 1'h0;
    end else begin
      _T_1534_3 <= _T_1534_2;
    end
    if (reset) begin
      _T_1546_0 <= 1'h0;
    end else begin
      _T_1546_0 <= _T_1367;
    end
    if (reset) begin
      _T_1546_1 <= 1'h0;
    end else begin
      _T_1546_1 <= _T_1546_0;
    end
    if (reset) begin
      _T_1546_2 <= 1'h0;
    end else begin
      _T_1546_2 <= _T_1546_1;
    end
    if (reset) begin
      _T_1546_3 <= 1'h0;
    end else begin
      _T_1546_3 <= _T_1546_2;
    end
    if (reset) begin
      _T_1558_0 <= 1'h0;
    end else begin
      _T_1558_0 <= _T_1465;
    end
    if (reset) begin
      _T_1558_1 <= 1'h0;
    end else begin
      _T_1558_1 <= _T_1558_0;
    end
    if (reset) begin
      _T_1558_2 <= 1'h0;
    end else begin
      _T_1558_2 <= _T_1558_1;
    end
    if (reset) begin
      _T_1558_3 <= 1'h0;
    end else begin
      _T_1558_3 <= _T_1558_2;
    end
    if (reset) begin
      _T_1570_0 <= 1'h0;
    end else begin
      _T_1570_0 <= _T_1563;
    end
    if (reset) begin
      _T_1570_1 <= 1'h0;
    end else begin
      _T_1570_1 <= _T_1570_0;
    end
    if (reset) begin
      _T_1570_2 <= 1'h0;
    end else begin
      _T_1570_2 <= _T_1570_1;
    end
    if (reset) begin
      _T_1570_3 <= 1'h0;
    end else begin
      _T_1570_3 <= _T_1570_2;
    end
    if (reset) begin
      _T_1585_0 <= 1'h0;
    end else begin
      _T_1585_0 <= _T_1580;
    end
    if (reset) begin
      _T_1585_1 <= 1'h0;
    end else begin
      _T_1585_1 <= _T_1585_0;
    end
    if (reset) begin
      _T_1585_2 <= 1'h0;
    end else begin
      _T_1585_2 <= _T_1585_1;
    end
    if (reset) begin
      _T_1594_0 <= 1'h0;
    end else begin
      _T_1594_0 <= _T_1589;
    end
    if (reset) begin
      _T_1594_1 <= 1'h0;
    end else begin
      _T_1594_1 <= _T_1594_0;
    end
    if (reset) begin
      _T_1594_2 <= 1'h0;
    end else begin
      _T_1594_2 <= _T_1594_1;
    end
    if (reset) begin
      _T_1603_0 <= 1'h0;
    end else begin
      _T_1603_0 <= _T_1598;
    end
    if (reset) begin
      _T_1603_1 <= 1'h0;
    end else begin
      _T_1603_1 <= _T_1603_0;
    end
    if (reset) begin
      _T_1603_2 <= 1'h0;
    end else begin
      _T_1603_2 <= _T_1603_1;
    end
    if (reset) begin
      _T_1612_0 <= 1'h0;
    end else begin
      _T_1612_0 <= _T_1607;
    end
    if (reset) begin
      _T_1612_1 <= 1'h0;
    end else begin
      _T_1612_1 <= _T_1612_0;
    end
    if (reset) begin
      _T_1612_2 <= 1'h0;
    end else begin
      _T_1612_2 <= _T_1612_1;
    end
    if (reset) begin
      _T_1621_0 <= 1'h0;
    end else begin
      _T_1621_0 <= _T_1616;
    end
    if (reset) begin
      _T_1621_1 <= 1'h0;
    end else begin
      _T_1621_1 <= _T_1621_0;
    end
    if (reset) begin
      _T_1621_2 <= 1'h0;
    end else begin
      _T_1621_2 <= _T_1621_1;
    end
    if (reset) begin
      _T_1630_0 <= 1'h0;
    end else begin
      _T_1630_0 <= _T_1625;
    end
    if (reset) begin
      _T_1630_1 <= 1'h0;
    end else begin
      _T_1630_1 <= _T_1630_0;
    end
    if (reset) begin
      _T_1630_2 <= 1'h0;
    end else begin
      _T_1630_2 <= _T_1630_1;
    end
    if (reset) begin
      _T_1639_0 <= 1'h0;
    end else begin
      _T_1639_0 <= _T_1634;
    end
    if (reset) begin
      _T_1639_1 <= 1'h0;
    end else begin
      _T_1639_1 <= _T_1639_0;
    end
    if (reset) begin
      _T_1639_2 <= 1'h0;
    end else begin
      _T_1639_2 <= _T_1639_1;
    end
    if (reset) begin
      _T_1648_0 <= 1'h0;
    end else begin
      _T_1648_0 <= _T_1643;
    end
    if (reset) begin
      _T_1648_1 <= 1'h0;
    end else begin
      _T_1648_1 <= _T_1648_0;
    end
    if (reset) begin
      _T_1648_2 <= 1'h0;
    end else begin
      _T_1648_2 <= _T_1648_1;
    end
    if (reset) begin
      _T_1657_0 <= 1'h0;
    end else begin
      _T_1657_0 <= _T_1652;
    end
    if (reset) begin
      _T_1657_1 <= 1'h0;
    end else begin
      _T_1657_1 <= _T_1657_0;
    end
    if (reset) begin
      _T_1657_2 <= 1'h0;
    end else begin
      _T_1657_2 <= _T_1657_1;
    end
    if (reset) begin
      _T_1666_0 <= 1'h0;
    end else begin
      _T_1666_0 <= _T_1661;
    end
    if (reset) begin
      _T_1666_1 <= 1'h0;
    end else begin
      _T_1666_1 <= _T_1666_0;
    end
    if (reset) begin
      _T_1666_2 <= 1'h0;
    end else begin
      _T_1666_2 <= _T_1666_1;
    end
    if (reset) begin
      _T_1675_0 <= 1'h0;
    end else begin
      _T_1675_0 <= _T_1670;
    end
    if (reset) begin
      _T_1675_1 <= 1'h0;
    end else begin
      _T_1675_1 <= _T_1675_0;
    end
    if (reset) begin
      _T_1675_2 <= 1'h0;
    end else begin
      _T_1675_2 <= _T_1675_1;
    end
    if (reset) begin
      _T_1684_0 <= 1'h0;
    end else begin
      _T_1684_0 <= _T_1679;
    end
    if (reset) begin
      _T_1684_1 <= 1'h0;
    end else begin
      _T_1684_1 <= _T_1684_0;
    end
    if (reset) begin
      _T_1684_2 <= 1'h0;
    end else begin
      _T_1684_2 <= _T_1684_1;
    end
    if (reset) begin
      _T_1693_0 <= 1'h0;
    end else begin
      _T_1693_0 <= _T_1688;
    end
    if (reset) begin
      _T_1693_1 <= 1'h0;
    end else begin
      _T_1693_1 <= _T_1693_0;
    end
    if (reset) begin
      _T_1693_2 <= 1'h0;
    end else begin
      _T_1693_2 <= _T_1693_1;
    end
    if (reset) begin
      _T_1702_0 <= 1'h0;
    end else begin
      _T_1702_0 <= _T_1697;
    end
    if (reset) begin
      _T_1702_1 <= 1'h0;
    end else begin
      _T_1702_1 <= _T_1702_0;
    end
    if (reset) begin
      _T_1702_2 <= 1'h0;
    end else begin
      _T_1702_2 <= _T_1702_1;
    end
    if (reset) begin
      _T_1711_0 <= 1'h0;
    end else begin
      _T_1711_0 <= _T_1706;
    end
    if (reset) begin
      _T_1711_1 <= 1'h0;
    end else begin
      _T_1711_1 <= _T_1711_0;
    end
    if (reset) begin
      _T_1711_2 <= 1'h0;
    end else begin
      _T_1711_2 <= _T_1711_1;
    end
    if (reset) begin
      _T_1720_0 <= 1'h0;
    end else begin
      _T_1720_0 <= _T_1715;
    end
    if (reset) begin
      _T_1720_1 <= 1'h0;
    end else begin
      _T_1720_1 <= _T_1720_0;
    end
    if (reset) begin
      _T_1720_2 <= 1'h0;
    end else begin
      _T_1720_2 <= _T_1720_1;
    end
    if (reset) begin
      _T_1722_0 <= 1'h0;
    end else begin
      _T_1722_0 <= io_exec_valid;
    end
    if (reset) begin
      _T_1722_1 <= 1'h0;
    end else begin
      _T_1722_1 <= _T_1722_0;
    end
    if (reset) begin
      _T_1722_2 <= 1'h0;
    end else begin
      _T_1722_2 <= _T_1722_1;
    end
    if (reset) begin
      _T_1722_3 <= 1'h0;
    end else begin
      _T_1722_3 <= _T_1722_2;
    end
    if (reset) begin
      _T_1722_4 <= 1'h0;
    end else begin
      _T_1722_4 <= _T_1722_3;
    end
    if (reset) begin
      _T_1722_5 <= 1'h0;
    end else begin
      _T_1722_5 <= _T_1722_4;
    end
    if (reset) begin
      _T_1722_6 <= 1'h0;
    end else begin
      _T_1722_6 <= _T_1722_5;
    end
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_1) begin
          $fwrite(32'h80000002,"exec_ctrl: Vec(%d, %d)\n",MultiDimTime_io_index_0,MultiDimTime_io_index_1); // @[pearray.scala 64:9]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_1) begin
          $fwrite(32'h80000002,"(%d, %d, %d, %d) ",PE_io_data_0_out_bits,PE_io_data_1_out_bits,PE_io_data_2_out_bits,PE_io_sig_stat2trans); // @[pearray.scala 170:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_1) begin
          $fwrite(32'h80000002,"(%d, %d, %d, %d) ",PE_1_io_data_0_out_bits,PE_1_io_data_1_out_bits,PE_1_io_data_2_out_bits,PE_1_io_sig_stat2trans); // @[pearray.scala 170:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_1) begin
          $fwrite(32'h80000002,"(%d, %d, %d, %d) ",PE_2_io_data_0_out_bits,PE_2_io_data_1_out_bits,PE_2_io_data_2_out_bits,PE_2_io_sig_stat2trans); // @[pearray.scala 170:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_1) begin
          $fwrite(32'h80000002,"(%d, %d, %d, %d) ",PE_3_io_data_0_out_bits,PE_3_io_data_1_out_bits,PE_3_io_data_2_out_bits,PE_3_io_sig_stat2trans); // @[pearray.scala 170:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_1) begin
          $fwrite(32'h80000002,"(%d, %d, %d, %d) ",PE_4_io_data_0_out_bits,PE_4_io_data_1_out_bits,PE_4_io_data_2_out_bits,PE_4_io_sig_stat2trans); // @[pearray.scala 170:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_1) begin
          $fwrite(32'h80000002,"(%d, %d, %d, %d) ",PE_5_io_data_0_out_bits,PE_5_io_data_1_out_bits,PE_5_io_data_2_out_bits,PE_5_io_sig_stat2trans); // @[pearray.scala 170:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_1) begin
          $fwrite(32'h80000002,"(%d, %d, %d, %d) ",PE_6_io_data_0_out_bits,PE_6_io_data_1_out_bits,PE_6_io_data_2_out_bits,PE_6_io_sig_stat2trans); // @[pearray.scala 170:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_1) begin
          $fwrite(32'h80000002,"(%d, %d, %d, %d) ",PE_7_io_data_0_out_bits,PE_7_io_data_1_out_bits,PE_7_io_data_2_out_bits,PE_7_io_sig_stat2trans); // @[pearray.scala 170:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_1) begin
          $fwrite(32'h80000002,"\n"); // @[pearray.scala 184:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_1) begin
          $fwrite(32'h80000002,"(%d, %d, %d, %d) ",PE_8_io_data_0_out_bits,PE_8_io_data_1_out_bits,PE_8_io_data_2_out_bits,PE_8_io_sig_stat2trans); // @[pearray.scala 170:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_1) begin
          $fwrite(32'h80000002,"(%d, %d, %d, %d) ",PE_9_io_data_0_out_bits,PE_9_io_data_1_out_bits,PE_9_io_data_2_out_bits,PE_9_io_sig_stat2trans); // @[pearray.scala 170:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_1) begin
          $fwrite(32'h80000002,"(%d, %d, %d, %d) ",PE_10_io_data_0_out_bits,PE_10_io_data_1_out_bits,PE_10_io_data_2_out_bits,PE_10_io_sig_stat2trans); // @[pearray.scala 170:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_1) begin
          $fwrite(32'h80000002,"(%d, %d, %d, %d) ",PE_11_io_data_0_out_bits,PE_11_io_data_1_out_bits,PE_11_io_data_2_out_bits,PE_11_io_sig_stat2trans); // @[pearray.scala 170:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_1) begin
          $fwrite(32'h80000002,"(%d, %d, %d, %d) ",PE_12_io_data_0_out_bits,PE_12_io_data_1_out_bits,PE_12_io_data_2_out_bits,PE_12_io_sig_stat2trans); // @[pearray.scala 170:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_1) begin
          $fwrite(32'h80000002,"(%d, %d, %d, %d) ",PE_13_io_data_0_out_bits,PE_13_io_data_1_out_bits,PE_13_io_data_2_out_bits,PE_13_io_sig_stat2trans); // @[pearray.scala 170:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_1) begin
          $fwrite(32'h80000002,"(%d, %d, %d, %d) ",PE_14_io_data_0_out_bits,PE_14_io_data_1_out_bits,PE_14_io_data_2_out_bits,PE_14_io_sig_stat2trans); // @[pearray.scala 170:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_1) begin
          $fwrite(32'h80000002,"(%d, %d, %d, %d) ",PE_15_io_data_0_out_bits,PE_15_io_data_1_out_bits,PE_15_io_data_2_out_bits,PE_15_io_sig_stat2trans); // @[pearray.scala 170:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_1) begin
          $fwrite(32'h80000002,"\n"); // @[pearray.scala 184:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_1) begin
          $fwrite(32'h80000002,"(%d, %d, %d, %d) ",PE_16_io_data_0_out_bits,PE_16_io_data_1_out_bits,PE_16_io_data_2_out_bits,PE_16_io_sig_stat2trans); // @[pearray.scala 170:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_1) begin
          $fwrite(32'h80000002,"(%d, %d, %d, %d) ",PE_17_io_data_0_out_bits,PE_17_io_data_1_out_bits,PE_17_io_data_2_out_bits,PE_17_io_sig_stat2trans); // @[pearray.scala 170:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_1) begin
          $fwrite(32'h80000002,"(%d, %d, %d, %d) ",PE_18_io_data_0_out_bits,PE_18_io_data_1_out_bits,PE_18_io_data_2_out_bits,PE_18_io_sig_stat2trans); // @[pearray.scala 170:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_1) begin
          $fwrite(32'h80000002,"(%d, %d, %d, %d) ",PE_19_io_data_0_out_bits,PE_19_io_data_1_out_bits,PE_19_io_data_2_out_bits,PE_19_io_sig_stat2trans); // @[pearray.scala 170:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_1) begin
          $fwrite(32'h80000002,"(%d, %d, %d, %d) ",PE_20_io_data_0_out_bits,PE_20_io_data_1_out_bits,PE_20_io_data_2_out_bits,PE_20_io_sig_stat2trans); // @[pearray.scala 170:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_1) begin
          $fwrite(32'h80000002,"(%d, %d, %d, %d) ",PE_21_io_data_0_out_bits,PE_21_io_data_1_out_bits,PE_21_io_data_2_out_bits,PE_21_io_sig_stat2trans); // @[pearray.scala 170:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_1) begin
          $fwrite(32'h80000002,"(%d, %d, %d, %d) ",PE_22_io_data_0_out_bits,PE_22_io_data_1_out_bits,PE_22_io_data_2_out_bits,PE_22_io_sig_stat2trans); // @[pearray.scala 170:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_1) begin
          $fwrite(32'h80000002,"(%d, %d, %d, %d) ",PE_23_io_data_0_out_bits,PE_23_io_data_1_out_bits,PE_23_io_data_2_out_bits,PE_23_io_sig_stat2trans); // @[pearray.scala 170:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_1) begin
          $fwrite(32'h80000002,"\n"); // @[pearray.scala 184:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_1) begin
          $fwrite(32'h80000002,"(%d, %d, %d, %d) ",PE_24_io_data_0_out_bits,PE_24_io_data_1_out_bits,PE_24_io_data_2_out_bits,PE_24_io_sig_stat2trans); // @[pearray.scala 170:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_1) begin
          $fwrite(32'h80000002,"(%d, %d, %d, %d) ",PE_25_io_data_0_out_bits,PE_25_io_data_1_out_bits,PE_25_io_data_2_out_bits,PE_25_io_sig_stat2trans); // @[pearray.scala 170:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_1) begin
          $fwrite(32'h80000002,"(%d, %d, %d, %d) ",PE_26_io_data_0_out_bits,PE_26_io_data_1_out_bits,PE_26_io_data_2_out_bits,PE_26_io_sig_stat2trans); // @[pearray.scala 170:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_1) begin
          $fwrite(32'h80000002,"(%d, %d, %d, %d) ",PE_27_io_data_0_out_bits,PE_27_io_data_1_out_bits,PE_27_io_data_2_out_bits,PE_27_io_sig_stat2trans); // @[pearray.scala 170:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_1) begin
          $fwrite(32'h80000002,"(%d, %d, %d, %d) ",PE_28_io_data_0_out_bits,PE_28_io_data_1_out_bits,PE_28_io_data_2_out_bits,PE_28_io_sig_stat2trans); // @[pearray.scala 170:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_1) begin
          $fwrite(32'h80000002,"(%d, %d, %d, %d) ",PE_29_io_data_0_out_bits,PE_29_io_data_1_out_bits,PE_29_io_data_2_out_bits,PE_29_io_sig_stat2trans); // @[pearray.scala 170:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_1) begin
          $fwrite(32'h80000002,"(%d, %d, %d, %d) ",PE_30_io_data_0_out_bits,PE_30_io_data_1_out_bits,PE_30_io_data_2_out_bits,PE_30_io_sig_stat2trans); // @[pearray.scala 170:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_1) begin
          $fwrite(32'h80000002,"(%d, %d, %d, %d) ",PE_31_io_data_0_out_bits,PE_31_io_data_1_out_bits,PE_31_io_data_2_out_bits,PE_31_io_sig_stat2trans); // @[pearray.scala 170:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_1) begin
          $fwrite(32'h80000002,"\n"); // @[pearray.scala 184:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_1) begin
          $fwrite(32'h80000002,"(%d, %d, %d, %d) ",PE_32_io_data_0_out_bits,PE_32_io_data_1_out_bits,PE_32_io_data_2_out_bits,PE_32_io_sig_stat2trans); // @[pearray.scala 170:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_1) begin
          $fwrite(32'h80000002,"(%d, %d, %d, %d) ",PE_33_io_data_0_out_bits,PE_33_io_data_1_out_bits,PE_33_io_data_2_out_bits,PE_33_io_sig_stat2trans); // @[pearray.scala 170:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_1) begin
          $fwrite(32'h80000002,"(%d, %d, %d, %d) ",PE_34_io_data_0_out_bits,PE_34_io_data_1_out_bits,PE_34_io_data_2_out_bits,PE_34_io_sig_stat2trans); // @[pearray.scala 170:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_1) begin
          $fwrite(32'h80000002,"(%d, %d, %d, %d) ",PE_35_io_data_0_out_bits,PE_35_io_data_1_out_bits,PE_35_io_data_2_out_bits,PE_35_io_sig_stat2trans); // @[pearray.scala 170:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_1) begin
          $fwrite(32'h80000002,"(%d, %d, %d, %d) ",PE_36_io_data_0_out_bits,PE_36_io_data_1_out_bits,PE_36_io_data_2_out_bits,PE_36_io_sig_stat2trans); // @[pearray.scala 170:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_1) begin
          $fwrite(32'h80000002,"(%d, %d, %d, %d) ",PE_37_io_data_0_out_bits,PE_37_io_data_1_out_bits,PE_37_io_data_2_out_bits,PE_37_io_sig_stat2trans); // @[pearray.scala 170:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_1) begin
          $fwrite(32'h80000002,"(%d, %d, %d, %d) ",PE_38_io_data_0_out_bits,PE_38_io_data_1_out_bits,PE_38_io_data_2_out_bits,PE_38_io_sig_stat2trans); // @[pearray.scala 170:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_1) begin
          $fwrite(32'h80000002,"(%d, %d, %d, %d) ",PE_39_io_data_0_out_bits,PE_39_io_data_1_out_bits,PE_39_io_data_2_out_bits,PE_39_io_sig_stat2trans); // @[pearray.scala 170:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_1) begin
          $fwrite(32'h80000002,"\n"); // @[pearray.scala 184:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_1) begin
          $fwrite(32'h80000002,"(%d, %d, %d, %d) ",PE_40_io_data_0_out_bits,PE_40_io_data_1_out_bits,PE_40_io_data_2_out_bits,PE_40_io_sig_stat2trans); // @[pearray.scala 170:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_1) begin
          $fwrite(32'h80000002,"(%d, %d, %d, %d) ",PE_41_io_data_0_out_bits,PE_41_io_data_1_out_bits,PE_41_io_data_2_out_bits,PE_41_io_sig_stat2trans); // @[pearray.scala 170:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_1) begin
          $fwrite(32'h80000002,"(%d, %d, %d, %d) ",PE_42_io_data_0_out_bits,PE_42_io_data_1_out_bits,PE_42_io_data_2_out_bits,PE_42_io_sig_stat2trans); // @[pearray.scala 170:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_1) begin
          $fwrite(32'h80000002,"(%d, %d, %d, %d) ",PE_43_io_data_0_out_bits,PE_43_io_data_1_out_bits,PE_43_io_data_2_out_bits,PE_43_io_sig_stat2trans); // @[pearray.scala 170:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_1) begin
          $fwrite(32'h80000002,"(%d, %d, %d, %d) ",PE_44_io_data_0_out_bits,PE_44_io_data_1_out_bits,PE_44_io_data_2_out_bits,PE_44_io_sig_stat2trans); // @[pearray.scala 170:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_1) begin
          $fwrite(32'h80000002,"(%d, %d, %d, %d) ",PE_45_io_data_0_out_bits,PE_45_io_data_1_out_bits,PE_45_io_data_2_out_bits,PE_45_io_sig_stat2trans); // @[pearray.scala 170:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_1) begin
          $fwrite(32'h80000002,"(%d, %d, %d, %d) ",PE_46_io_data_0_out_bits,PE_46_io_data_1_out_bits,PE_46_io_data_2_out_bits,PE_46_io_sig_stat2trans); // @[pearray.scala 170:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_1) begin
          $fwrite(32'h80000002,"(%d, %d, %d, %d) ",PE_47_io_data_0_out_bits,PE_47_io_data_1_out_bits,PE_47_io_data_2_out_bits,PE_47_io_sig_stat2trans); // @[pearray.scala 170:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_1) begin
          $fwrite(32'h80000002,"\n"); // @[pearray.scala 184:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_1) begin
          $fwrite(32'h80000002,"(%d, %d, %d, %d) ",PE_48_io_data_0_out_bits,PE_48_io_data_1_out_bits,PE_48_io_data_2_out_bits,PE_48_io_sig_stat2trans); // @[pearray.scala 170:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_1) begin
          $fwrite(32'h80000002,"(%d, %d, %d, %d) ",PE_49_io_data_0_out_bits,PE_49_io_data_1_out_bits,PE_49_io_data_2_out_bits,PE_49_io_sig_stat2trans); // @[pearray.scala 170:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_1) begin
          $fwrite(32'h80000002,"(%d, %d, %d, %d) ",PE_50_io_data_0_out_bits,PE_50_io_data_1_out_bits,PE_50_io_data_2_out_bits,PE_50_io_sig_stat2trans); // @[pearray.scala 170:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_1) begin
          $fwrite(32'h80000002,"(%d, %d, %d, %d) ",PE_51_io_data_0_out_bits,PE_51_io_data_1_out_bits,PE_51_io_data_2_out_bits,PE_51_io_sig_stat2trans); // @[pearray.scala 170:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_1) begin
          $fwrite(32'h80000002,"(%d, %d, %d, %d) ",PE_52_io_data_0_out_bits,PE_52_io_data_1_out_bits,PE_52_io_data_2_out_bits,PE_52_io_sig_stat2trans); // @[pearray.scala 170:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_1) begin
          $fwrite(32'h80000002,"(%d, %d, %d, %d) ",PE_53_io_data_0_out_bits,PE_53_io_data_1_out_bits,PE_53_io_data_2_out_bits,PE_53_io_sig_stat2trans); // @[pearray.scala 170:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_1) begin
          $fwrite(32'h80000002,"(%d, %d, %d, %d) ",PE_54_io_data_0_out_bits,PE_54_io_data_1_out_bits,PE_54_io_data_2_out_bits,PE_54_io_sig_stat2trans); // @[pearray.scala 170:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_1) begin
          $fwrite(32'h80000002,"(%d, %d, %d, %d) ",PE_55_io_data_0_out_bits,PE_55_io_data_1_out_bits,PE_55_io_data_2_out_bits,PE_55_io_sig_stat2trans); // @[pearray.scala 170:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_1) begin
          $fwrite(32'h80000002,"\n"); // @[pearray.scala 184:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_1) begin
          $fwrite(32'h80000002,"(%d, %d, %d, %d) ",PE_56_io_data_0_out_bits,PE_56_io_data_1_out_bits,PE_56_io_data_2_out_bits,PE_56_io_sig_stat2trans); // @[pearray.scala 170:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_1) begin
          $fwrite(32'h80000002,"(%d, %d, %d, %d) ",PE_57_io_data_0_out_bits,PE_57_io_data_1_out_bits,PE_57_io_data_2_out_bits,PE_57_io_sig_stat2trans); // @[pearray.scala 170:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_1) begin
          $fwrite(32'h80000002,"(%d, %d, %d, %d) ",PE_58_io_data_0_out_bits,PE_58_io_data_1_out_bits,PE_58_io_data_2_out_bits,PE_58_io_sig_stat2trans); // @[pearray.scala 170:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_1) begin
          $fwrite(32'h80000002,"(%d, %d, %d, %d) ",PE_59_io_data_0_out_bits,PE_59_io_data_1_out_bits,PE_59_io_data_2_out_bits,PE_59_io_sig_stat2trans); // @[pearray.scala 170:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_1) begin
          $fwrite(32'h80000002,"(%d, %d, %d, %d) ",PE_60_io_data_0_out_bits,PE_60_io_data_1_out_bits,PE_60_io_data_2_out_bits,PE_60_io_sig_stat2trans); // @[pearray.scala 170:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_1) begin
          $fwrite(32'h80000002,"(%d, %d, %d, %d) ",PE_61_io_data_0_out_bits,PE_61_io_data_1_out_bits,PE_61_io_data_2_out_bits,PE_61_io_sig_stat2trans); // @[pearray.scala 170:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_1) begin
          $fwrite(32'h80000002,"(%d, %d, %d, %d) ",PE_62_io_data_0_out_bits,PE_62_io_data_1_out_bits,PE_62_io_data_2_out_bits,PE_62_io_sig_stat2trans); // @[pearray.scala 170:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_1) begin
          $fwrite(32'h80000002,"(%d, %d, %d, %d) ",PE_63_io_data_0_out_bits,PE_63_io_data_1_out_bits,PE_63_io_data_2_out_bits,PE_63_io_sig_stat2trans); // @[pearray.scala 170:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_1) begin
          $fwrite(32'h80000002,"\n"); // @[pearray.scala 184:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_1) begin
          $fwrite(32'h80000002,"(%d, %d, %d, %d) ",PE_64_io_data_0_out_bits,PE_64_io_data_1_out_bits,PE_64_io_data_2_out_bits,PE_64_io_sig_stat2trans); // @[pearray.scala 170:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_1) begin
          $fwrite(32'h80000002,"(%d, %d, %d, %d) ",PE_65_io_data_0_out_bits,PE_65_io_data_1_out_bits,PE_65_io_data_2_out_bits,PE_65_io_sig_stat2trans); // @[pearray.scala 170:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_1) begin
          $fwrite(32'h80000002,"(%d, %d, %d, %d) ",PE_66_io_data_0_out_bits,PE_66_io_data_1_out_bits,PE_66_io_data_2_out_bits,PE_66_io_sig_stat2trans); // @[pearray.scala 170:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_1) begin
          $fwrite(32'h80000002,"(%d, %d, %d, %d) ",PE_67_io_data_0_out_bits,PE_67_io_data_1_out_bits,PE_67_io_data_2_out_bits,PE_67_io_sig_stat2trans); // @[pearray.scala 170:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_1) begin
          $fwrite(32'h80000002,"(%d, %d, %d, %d) ",PE_68_io_data_0_out_bits,PE_68_io_data_1_out_bits,PE_68_io_data_2_out_bits,PE_68_io_sig_stat2trans); // @[pearray.scala 170:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_1) begin
          $fwrite(32'h80000002,"(%d, %d, %d, %d) ",PE_69_io_data_0_out_bits,PE_69_io_data_1_out_bits,PE_69_io_data_2_out_bits,PE_69_io_sig_stat2trans); // @[pearray.scala 170:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_1) begin
          $fwrite(32'h80000002,"(%d, %d, %d, %d) ",PE_70_io_data_0_out_bits,PE_70_io_data_1_out_bits,PE_70_io_data_2_out_bits,PE_70_io_sig_stat2trans); // @[pearray.scala 170:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_1) begin
          $fwrite(32'h80000002,"(%d, %d, %d, %d) ",PE_71_io_data_0_out_bits,PE_71_io_data_1_out_bits,PE_71_io_data_2_out_bits,PE_71_io_sig_stat2trans); // @[pearray.scala 170:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_1) begin
          $fwrite(32'h80000002,"\n"); // @[pearray.scala 184:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_1) begin
          $fwrite(32'h80000002,"(%d, %d, %d, %d) ",PE_72_io_data_0_out_bits,PE_72_io_data_1_out_bits,PE_72_io_data_2_out_bits,PE_72_io_sig_stat2trans); // @[pearray.scala 170:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_1) begin
          $fwrite(32'h80000002,"(%d, %d, %d, %d) ",PE_73_io_data_0_out_bits,PE_73_io_data_1_out_bits,PE_73_io_data_2_out_bits,PE_73_io_sig_stat2trans); // @[pearray.scala 170:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_1) begin
          $fwrite(32'h80000002,"(%d, %d, %d, %d) ",PE_74_io_data_0_out_bits,PE_74_io_data_1_out_bits,PE_74_io_data_2_out_bits,PE_74_io_sig_stat2trans); // @[pearray.scala 170:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_1) begin
          $fwrite(32'h80000002,"(%d, %d, %d, %d) ",PE_75_io_data_0_out_bits,PE_75_io_data_1_out_bits,PE_75_io_data_2_out_bits,PE_75_io_sig_stat2trans); // @[pearray.scala 170:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_1) begin
          $fwrite(32'h80000002,"(%d, %d, %d, %d) ",PE_76_io_data_0_out_bits,PE_76_io_data_1_out_bits,PE_76_io_data_2_out_bits,PE_76_io_sig_stat2trans); // @[pearray.scala 170:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_1) begin
          $fwrite(32'h80000002,"(%d, %d, %d, %d) ",PE_77_io_data_0_out_bits,PE_77_io_data_1_out_bits,PE_77_io_data_2_out_bits,PE_77_io_sig_stat2trans); // @[pearray.scala 170:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_1) begin
          $fwrite(32'h80000002,"(%d, %d, %d, %d) ",PE_78_io_data_0_out_bits,PE_78_io_data_1_out_bits,PE_78_io_data_2_out_bits,PE_78_io_sig_stat2trans); // @[pearray.scala 170:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_1) begin
          $fwrite(32'h80000002,"(%d, %d, %d, %d) ",PE_79_io_data_0_out_bits,PE_79_io_data_1_out_bits,PE_79_io_data_2_out_bits,PE_79_io_sig_stat2trans); // @[pearray.scala 170:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_1) begin
          $fwrite(32'h80000002,"\n"); // @[pearray.scala 184:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_1) begin
          $fwrite(32'h80000002,"(%d, %d, %d, %d) ",PE_80_io_data_0_out_bits,PE_80_io_data_1_out_bits,PE_80_io_data_2_out_bits,PE_80_io_sig_stat2trans); // @[pearray.scala 170:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_1) begin
          $fwrite(32'h80000002,"(%d, %d, %d, %d) ",PE_81_io_data_0_out_bits,PE_81_io_data_1_out_bits,PE_81_io_data_2_out_bits,PE_81_io_sig_stat2trans); // @[pearray.scala 170:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_1) begin
          $fwrite(32'h80000002,"(%d, %d, %d, %d) ",PE_82_io_data_0_out_bits,PE_82_io_data_1_out_bits,PE_82_io_data_2_out_bits,PE_82_io_sig_stat2trans); // @[pearray.scala 170:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_1) begin
          $fwrite(32'h80000002,"(%d, %d, %d, %d) ",PE_83_io_data_0_out_bits,PE_83_io_data_1_out_bits,PE_83_io_data_2_out_bits,PE_83_io_sig_stat2trans); // @[pearray.scala 170:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_1) begin
          $fwrite(32'h80000002,"(%d, %d, %d, %d) ",PE_84_io_data_0_out_bits,PE_84_io_data_1_out_bits,PE_84_io_data_2_out_bits,PE_84_io_sig_stat2trans); // @[pearray.scala 170:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_1) begin
          $fwrite(32'h80000002,"(%d, %d, %d, %d) ",PE_85_io_data_0_out_bits,PE_85_io_data_1_out_bits,PE_85_io_data_2_out_bits,PE_85_io_sig_stat2trans); // @[pearray.scala 170:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_1) begin
          $fwrite(32'h80000002,"(%d, %d, %d, %d) ",PE_86_io_data_0_out_bits,PE_86_io_data_1_out_bits,PE_86_io_data_2_out_bits,PE_86_io_sig_stat2trans); // @[pearray.scala 170:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_1) begin
          $fwrite(32'h80000002,"(%d, %d, %d, %d) ",PE_87_io_data_0_out_bits,PE_87_io_data_1_out_bits,PE_87_io_data_2_out_bits,PE_87_io_sig_stat2trans); // @[pearray.scala 170:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_1) begin
          $fwrite(32'h80000002,"\n"); // @[pearray.scala 184:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_1) begin
          $fwrite(32'h80000002,"(%d, %d, %d, %d) ",PE_88_io_data_0_out_bits,PE_88_io_data_1_out_bits,PE_88_io_data_2_out_bits,PE_88_io_sig_stat2trans); // @[pearray.scala 170:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_1) begin
          $fwrite(32'h80000002,"(%d, %d, %d, %d) ",PE_89_io_data_0_out_bits,PE_89_io_data_1_out_bits,PE_89_io_data_2_out_bits,PE_89_io_sig_stat2trans); // @[pearray.scala 170:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_1) begin
          $fwrite(32'h80000002,"(%d, %d, %d, %d) ",PE_90_io_data_0_out_bits,PE_90_io_data_1_out_bits,PE_90_io_data_2_out_bits,PE_90_io_sig_stat2trans); // @[pearray.scala 170:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_1) begin
          $fwrite(32'h80000002,"(%d, %d, %d, %d) ",PE_91_io_data_0_out_bits,PE_91_io_data_1_out_bits,PE_91_io_data_2_out_bits,PE_91_io_sig_stat2trans); // @[pearray.scala 170:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_1) begin
          $fwrite(32'h80000002,"(%d, %d, %d, %d) ",PE_92_io_data_0_out_bits,PE_92_io_data_1_out_bits,PE_92_io_data_2_out_bits,PE_92_io_sig_stat2trans); // @[pearray.scala 170:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_1) begin
          $fwrite(32'h80000002,"(%d, %d, %d, %d) ",PE_93_io_data_0_out_bits,PE_93_io_data_1_out_bits,PE_93_io_data_2_out_bits,PE_93_io_sig_stat2trans); // @[pearray.scala 170:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_1) begin
          $fwrite(32'h80000002,"(%d, %d, %d, %d) ",PE_94_io_data_0_out_bits,PE_94_io_data_1_out_bits,PE_94_io_data_2_out_bits,PE_94_io_sig_stat2trans); // @[pearray.scala 170:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_1) begin
          $fwrite(32'h80000002,"(%d, %d, %d, %d) ",PE_95_io_data_0_out_bits,PE_95_io_data_1_out_bits,PE_95_io_data_2_out_bits,PE_95_io_sig_stat2trans); // @[pearray.scala 170:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_1) begin
          $fwrite(32'h80000002,"\n"); // @[pearray.scala 184:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_1) begin
          $fwrite(32'h80000002,"(%d, %d, %d, %d) ",PE_96_io_data_0_out_bits,PE_96_io_data_1_out_bits,PE_96_io_data_2_out_bits,PE_96_io_sig_stat2trans); // @[pearray.scala 170:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_1) begin
          $fwrite(32'h80000002,"(%d, %d, %d, %d) ",PE_97_io_data_0_out_bits,PE_97_io_data_1_out_bits,PE_97_io_data_2_out_bits,PE_97_io_sig_stat2trans); // @[pearray.scala 170:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_1) begin
          $fwrite(32'h80000002,"(%d, %d, %d, %d) ",PE_98_io_data_0_out_bits,PE_98_io_data_1_out_bits,PE_98_io_data_2_out_bits,PE_98_io_sig_stat2trans); // @[pearray.scala 170:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_1) begin
          $fwrite(32'h80000002,"(%d, %d, %d, %d) ",PE_99_io_data_0_out_bits,PE_99_io_data_1_out_bits,PE_99_io_data_2_out_bits,PE_99_io_sig_stat2trans); // @[pearray.scala 170:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_1) begin
          $fwrite(32'h80000002,"(%d, %d, %d, %d) ",PE_100_io_data_0_out_bits,PE_100_io_data_1_out_bits,PE_100_io_data_2_out_bits,PE_100_io_sig_stat2trans); // @[pearray.scala 170:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_1) begin
          $fwrite(32'h80000002,"(%d, %d, %d, %d) ",PE_101_io_data_0_out_bits,PE_101_io_data_1_out_bits,PE_101_io_data_2_out_bits,PE_101_io_sig_stat2trans); // @[pearray.scala 170:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_1) begin
          $fwrite(32'h80000002,"(%d, %d, %d, %d) ",PE_102_io_data_0_out_bits,PE_102_io_data_1_out_bits,PE_102_io_data_2_out_bits,PE_102_io_sig_stat2trans); // @[pearray.scala 170:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_1) begin
          $fwrite(32'h80000002,"(%d, %d, %d, %d) ",PE_103_io_data_0_out_bits,PE_103_io_data_1_out_bits,PE_103_io_data_2_out_bits,PE_103_io_sig_stat2trans); // @[pearray.scala 170:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_1) begin
          $fwrite(32'h80000002,"\n"); // @[pearray.scala 184:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_1) begin
          $fwrite(32'h80000002,"(%d, %d, %d, %d) ",PE_104_io_data_0_out_bits,PE_104_io_data_1_out_bits,PE_104_io_data_2_out_bits,PE_104_io_sig_stat2trans); // @[pearray.scala 170:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_1) begin
          $fwrite(32'h80000002,"(%d, %d, %d, %d) ",PE_105_io_data_0_out_bits,PE_105_io_data_1_out_bits,PE_105_io_data_2_out_bits,PE_105_io_sig_stat2trans); // @[pearray.scala 170:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_1) begin
          $fwrite(32'h80000002,"(%d, %d, %d, %d) ",PE_106_io_data_0_out_bits,PE_106_io_data_1_out_bits,PE_106_io_data_2_out_bits,PE_106_io_sig_stat2trans); // @[pearray.scala 170:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_1) begin
          $fwrite(32'h80000002,"(%d, %d, %d, %d) ",PE_107_io_data_0_out_bits,PE_107_io_data_1_out_bits,PE_107_io_data_2_out_bits,PE_107_io_sig_stat2trans); // @[pearray.scala 170:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_1) begin
          $fwrite(32'h80000002,"(%d, %d, %d, %d) ",PE_108_io_data_0_out_bits,PE_108_io_data_1_out_bits,PE_108_io_data_2_out_bits,PE_108_io_sig_stat2trans); // @[pearray.scala 170:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_1) begin
          $fwrite(32'h80000002,"(%d, %d, %d, %d) ",PE_109_io_data_0_out_bits,PE_109_io_data_1_out_bits,PE_109_io_data_2_out_bits,PE_109_io_sig_stat2trans); // @[pearray.scala 170:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_1) begin
          $fwrite(32'h80000002,"(%d, %d, %d, %d) ",PE_110_io_data_0_out_bits,PE_110_io_data_1_out_bits,PE_110_io_data_2_out_bits,PE_110_io_sig_stat2trans); // @[pearray.scala 170:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_1) begin
          $fwrite(32'h80000002,"(%d, %d, %d, %d) ",PE_111_io_data_0_out_bits,PE_111_io_data_1_out_bits,PE_111_io_data_2_out_bits,PE_111_io_sig_stat2trans); // @[pearray.scala 170:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_1) begin
          $fwrite(32'h80000002,"\n"); // @[pearray.scala 184:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_1) begin
          $fwrite(32'h80000002,"(%d, %d, %d, %d) ",PE_112_io_data_0_out_bits,PE_112_io_data_1_out_bits,PE_112_io_data_2_out_bits,PE_112_io_sig_stat2trans); // @[pearray.scala 170:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_1) begin
          $fwrite(32'h80000002,"(%d, %d, %d, %d) ",PE_113_io_data_0_out_bits,PE_113_io_data_1_out_bits,PE_113_io_data_2_out_bits,PE_113_io_sig_stat2trans); // @[pearray.scala 170:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_1) begin
          $fwrite(32'h80000002,"(%d, %d, %d, %d) ",PE_114_io_data_0_out_bits,PE_114_io_data_1_out_bits,PE_114_io_data_2_out_bits,PE_114_io_sig_stat2trans); // @[pearray.scala 170:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_1) begin
          $fwrite(32'h80000002,"(%d, %d, %d, %d) ",PE_115_io_data_0_out_bits,PE_115_io_data_1_out_bits,PE_115_io_data_2_out_bits,PE_115_io_sig_stat2trans); // @[pearray.scala 170:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_1) begin
          $fwrite(32'h80000002,"(%d, %d, %d, %d) ",PE_116_io_data_0_out_bits,PE_116_io_data_1_out_bits,PE_116_io_data_2_out_bits,PE_116_io_sig_stat2trans); // @[pearray.scala 170:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_1) begin
          $fwrite(32'h80000002,"(%d, %d, %d, %d) ",PE_117_io_data_0_out_bits,PE_117_io_data_1_out_bits,PE_117_io_data_2_out_bits,PE_117_io_sig_stat2trans); // @[pearray.scala 170:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_1) begin
          $fwrite(32'h80000002,"(%d, %d, %d, %d) ",PE_118_io_data_0_out_bits,PE_118_io_data_1_out_bits,PE_118_io_data_2_out_bits,PE_118_io_sig_stat2trans); // @[pearray.scala 170:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_1) begin
          $fwrite(32'h80000002,"(%d, %d, %d, %d) ",PE_119_io_data_0_out_bits,PE_119_io_data_1_out_bits,PE_119_io_data_2_out_bits,PE_119_io_sig_stat2trans); // @[pearray.scala 170:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_1) begin
          $fwrite(32'h80000002,"\n"); // @[pearray.scala 184:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_1) begin
          $fwrite(32'h80000002,"(%d, %d, %d, %d) ",PE_120_io_data_0_out_bits,PE_120_io_data_1_out_bits,PE_120_io_data_2_out_bits,PE_120_io_sig_stat2trans); // @[pearray.scala 170:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_1) begin
          $fwrite(32'h80000002,"(%d, %d, %d, %d) ",PE_121_io_data_0_out_bits,PE_121_io_data_1_out_bits,PE_121_io_data_2_out_bits,PE_121_io_sig_stat2trans); // @[pearray.scala 170:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_1) begin
          $fwrite(32'h80000002,"(%d, %d, %d, %d) ",PE_122_io_data_0_out_bits,PE_122_io_data_1_out_bits,PE_122_io_data_2_out_bits,PE_122_io_sig_stat2trans); // @[pearray.scala 170:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_1) begin
          $fwrite(32'h80000002,"(%d, %d, %d, %d) ",PE_123_io_data_0_out_bits,PE_123_io_data_1_out_bits,PE_123_io_data_2_out_bits,PE_123_io_sig_stat2trans); // @[pearray.scala 170:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_1) begin
          $fwrite(32'h80000002,"(%d, %d, %d, %d) ",PE_124_io_data_0_out_bits,PE_124_io_data_1_out_bits,PE_124_io_data_2_out_bits,PE_124_io_sig_stat2trans); // @[pearray.scala 170:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_1) begin
          $fwrite(32'h80000002,"(%d, %d, %d, %d) ",PE_125_io_data_0_out_bits,PE_125_io_data_1_out_bits,PE_125_io_data_2_out_bits,PE_125_io_sig_stat2trans); // @[pearray.scala 170:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_1) begin
          $fwrite(32'h80000002,"(%d, %d, %d, %d) ",PE_126_io_data_0_out_bits,PE_126_io_data_1_out_bits,PE_126_io_data_2_out_bits,PE_126_io_sig_stat2trans); // @[pearray.scala 170:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_1) begin
          $fwrite(32'h80000002,"(%d, %d, %d, %d) ",PE_127_io_data_0_out_bits,PE_127_io_data_1_out_bits,PE_127_io_data_2_out_bits,PE_127_io_sig_stat2trans); // @[pearray.scala 170:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_1) begin
          $fwrite(32'h80000002,"\n"); // @[pearray.scala 184:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
  end
endmodule
